`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
TUg3INHh1m7IhzJTWhl4hakhjur7Vc43ogrhEddqQLKQ5cTmQJLyY/O39MHvxAMR2gKZYkMnwG2l
6cfBg6sy6w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Y/ia27A6wO8jmiJeDD7eisp/o0DINS9aBVInHA54TUKf2WoIq6hh9BVkHnKwsRC6y0ISNQHYfAzE
PTfro7nWLiogO1UdUR6Fdg0dugY297GMGNSgJp4hSjDcncspoXCIzLXdW36IFe/bIH2I6rVCdQGq
Bfb5Gy8ISAcPnQqsvfA=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
kz0wef7kcYmKk02nW3FHEht391vWQJY92Du/ZIt2m7OdokLfO6Gv5DKbZwOuyO+yXdcUUdWHG1Hg
t7gRWxEAkdlL4/9TviviX6GS9QtH9m8xJMYQY/3evLZuJv2spaJpj9XdTT9hQlWB3KOO/c4zrwkZ
4xmqwjxejGJsb+FM5sQ=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dkOPiv2V30YAr2yuyXphkE0lv+yYw3tHqA0yhJuJHSglEGmP0QTtSBhDMb+PGYV8NkSI8H4eVQnW
syXqKR2vhzWnJ0zRCtYlN/vMwjrZm35SHeCGC3CWsCXPg5fWlXJzxzDU4vP5OD4maGH8Ec1mMktz
gRtGcXleZSmjeO8rz4N7Zl+e7irHttUbvM4i2n84/VDlVWomp1+ZWh9VIiNadiVaF4GeyDmNDujq
KQ5joBbbe4y2hoQTmu/mtfDUMZGGvUoImw+vazPIlVHH7z5MXdEpWiEKnH14qDniwjKNjq35y1au
oZwXSsG5YkjKitE/OpWH3/uszWGUyrd02WCk7g==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YPeWnh+rwbGP5pImDI2d2//p4f/IpBCUCuKd/hCDk+2PHES852iLZdoJloFPd1161LDanxCbRI/P
1nJbZi1obBy3B4ujpRc/a43DfJ7dxQHZtNjYKs9a//VCBS+23vBkqK8aImNg1Enfw1pvrz0j2FHW
6mOF4jYRiH5WXOIIuBHFpcloerzd0g9AWQUxk/T+WCSCqmYWUEWg517jiOu9LvsqInAOCZ5t0SWx
1A5jeWyL+aVl7ZT62sEEoT6kmD5KQH/kGkUI9nUWAJWa2/k8yR8JxLoz3s/KFTMxpyrcHKw2Mba6
kP0rB/IanjAxmkWkkMe1p+USCoEpuIy40jLfFA==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2015_12", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RAvb/4vlo/jbWHAYh5QgcKvlffxbz7XViXDEv3yRgfG8bjy/C4S5r75Las5nWMxVHPrwZeDhcP3y
eWa+WDaWFUlrAa+9O9M4rBFwyH6vPJbUtAoKNZ7YapE5ME95Y4BKJQml4a6fc9hGkDkuDTohQL+e
h1h5j2N9YkWtTKH92l+ACHoeTq3jJ7tMmqXWKNWTJN+Wsc2eZhJhClQDjPMSNa3YztWgvs7raemX
fIP1EibAwQWW24hS/XYADD61gRmAHEtBDkKgnD8twsgno/WaAeXts9/ZgPRMk/yeorVQWfEagZMk
7092cD8GLSfd1pkbwQlcvmGKY4sXaCSxbhTWwA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 126032)
`protect data_block
3xwWy/6MRkRZeShS+gzVnyCgu6hmxBCku8OmzHxtEmPfQhdBrJUFZbsyilcsmXF9fxe07WZOuEfd
29eDCusqS6+GDkQa1fObrFpDTlGsg/zuZPKlOxbgj2ogFnMxnIt9mTUOm/CSQZjfBQ7ygkuzC+46
LvVkp2t9HZAvuSAyMZznF4cqG5AAhJvQU1qqZfPY0AR7DCBAQy31VXzjIVWQ26+QZ0TGIhk1ERrN
IJFDiUlNRrtxLq9WMMPF9Oy2fUuKxCbahSnogmQZTAWUYCja/VXw0bqyhlD4MXbIHXTM3X+aBCe/
5QSNpZFK3LtLbQe68WvdwSyURbOkc2SzWP/a6odnSOay98eYKLf7Zq6mEXmWGJTlFH5lDdsIO94e
S3v5LZIAnPAG7jPY1Ljr66SrMRz1EPDbrfQAvu6rmkTEAqvreWAFHrJhAshRav7gbDA1MZ981/xB
b6kEszqjckJogNAa6Xl5kJurk7cpJABroH2dFytHhVy4ze/+fwesoHFV/Q3HZiAHFKEM9DtpLo2s
qTltHTlgUzI6hS09RD6/zKLs6TcGgfgAR71IUe0mpuvr/pF90dBzgyIMr0ujtTjunzOLeOAeChWk
RBxBgjAiFk5KsOeGA0jtyegJ5UN0Ol0JUlRmNCzL6kiajDqOsdvqZSN5ni8eUtnUy8W4Afkerlxz
CmBiC/d1aBqVPxN5ppWmZEGvQWjujgx6gf1dj13x77Af7FfZOs9WqVRhSJJrWMO4fJQpXbUMoZSz
Xq3bD3IlXclwTu4LkrwFD6EKQMdViPgZqIhu3ppfS3yQhn+g1GbhN7Hc9wgNYmm3XDOXH3wzV531
8LoBGd3Msr7am/v9mOeNGt6Xx4z5I7RPDkffQFOGsoprm4vCHMzurHlYzWHPUdDqDvJ7+b54Z5C8
DaxyLh+lLT9+/lDs4h+qH7yfL3eeqZBN2zDjrwjvlsnsIMnyVQgOPFC1dUYwkm88Vah6G7O0NuH0
UYdBDwSqdGyqnS6eHsB4ia+Y23Qd75J5twb9/lQGl0dr8fPaBdpxfZmq9LGRpdrBmvzngwEzR48T
MxBVge0eDEnAaFnCNAI3AUE3mm34o9aH7piZNAA9b+JO7SAArLNZ6wgl2717AGAZ3TpU4bfmxVot
7Y6R7h23pTrqVY44GJdgKRBQ6DQ2SPnCwQRi4Q5/XPZDCKkr8gz1aseDxAtFQxdayMOHeQ9kCcp+
gQ2PoxKwDSVg8z3QjRFTvWFlohpIowOw2pZl7wU5RVRSPAXYGKYq+RjvRgrQAvIvxVOBrnHH11TO
826DmNQ3gbHIys2Y2kpesvU1cbackMog70cOelnYP/my6ZtOKRPwCwTeKNAPFmJgLwhWxmhKY8I9
xG/+ztD9I8FHWqozE3cxG1qhNPTT+dZ2x0S9fFA/INZnGGv0j1Em6zp6sKLTQIghWfde1SaTz+qK
eOY5fU6Tgm4sIoV4nkz6LLRe8euzFyguFKDmFb2dH5hHk/oqGVB7+76y79TBfSFu00Ck9BPaB3hK
oMvRy5+CE0/zGYz39+Z0gbBK5/YVJZ6Yx7BKlG5GKtj9fOjUCbJbPqgFqoAJFsJvBRCTalwWIwxi
+47WnMnGA0mvSei/b16TrBI0d4nBMP4ydy5bNkSpUZNhfh17j+2DMhCpnsgvPTLMBM7qwLwbaSF4
Jl5U7eub2uJlvGDWM3j4icIkr2bfcnrhrLxF0sx06oz7jtjIBnME/CQaKU8GshBpQjLypwgIlT3w
DWhKSRxRMHqq4Gi9QqXJBBIUWtiq8ziqfRGyHZkTT6c/Vjw4/gTWZ79eYQQ01+DVjp7RzA9KfLBT
ld8tHNOQPwd2+gSGnp8zXhb2t4r4M6ujH6IMPIWgcWGmygzc1MhNRH19w7ysRu8rEXVkEhwG8Pb9
W4HICsubX8/PId9YvwsXYImeIW0wdUNSbZTxIIkfK55Go0NYXSrT0ap4CEPWzA7ZdWu8VJshAilj
l+xM7KfsSNECpCRrBjG0RQrWsPMbH1B7E7IALtEFRjztXZzL9/7/+e4gGbIz5pfLybmeqqGhKzIR
UH6Tlxm/8X77Km0ksofduOB/QyLZ6+FnjIFJ5GdzLairynMIW89p3LJO9YcOCX3Z4QqzOQdCn37L
z8w0VxkfKeyKdTvcErn66yYcbV/9MFs/WL95UYAVYQOCw04b5992lULw3F5DVxkd5AwnfY0bE9RQ
U1HEAOxgNpz+Qh2ipGvsDyRPyfW91WhnS/DmawyYbuP3FSm4r2knmPbd/U2TPkTlSFnItpl0ltZ9
iFepSSPjiXv2ZO1JWPcBt7LMYq8iR4geb3xR5WbpIAqb+LXu0dhsJP1SxqHSkdKfVAPHCK2nyyWy
J8lO0B7zAUNvXnC+OUmGy60Rt0WC/2IaQv3dt/He/lGxndUaiFzFK6M+JAWOJx4GOi96Lf0DpiJY
+3NdKiXELwi/GNpIRZilW/pJwmB5SLnksI9Nbb1S0Jem8zKUHRQrCA+qgGfO390iELI+AByRh5HJ
vynXaQssjmt6zbe07zyrc8UwLNaud6BojgjT7wKq5oKCHVHfv70W4oqVeXyH1liz7knBRX3iPsFI
GXqKwk7D+UYUx9f08715lPWRf9oMZxTsVGgWVdnECG5kPSp0tGZKK2h8PS+hgnCcE4y2aFoyfQlA
wb4z1zQf2wKd89dDx0Zqup2btvzgY5U20sn+zzZocHMVYn/b9Mb8HkdiyVC4urvaxksPYhiJB+R4
xtceUdEWH07u2hnhoUJCQ7cBwH05NAQDwELAH37SWosxSTi4X7sJ5/lxIbHvD8Izwv8/iwrYlXPh
hGilVMxUOjWQGI5LpjYFzwX/qsSCY3feFwnIVdZN5k8Ip/LwyuvywrI18nmfrqnxBgwczK661RJx
sxg541vHBZHlYIkSaBOEte224IOSmurKEhPYSRzWBvD2CELtIKpFVj+okmUYgYH3grOrHdE9NXTV
C0Asqzec2j6p44zM7VN+mpxrqapFfw2VQOcqx/qlrZ5nP1HvHi6P7xikvFsPUnnJWqf20F2x/Qul
HHM0wNIsvyxcy/+Fi4TBVjpe7mv+LD5ajwNr66IAS6Cb1y3FfB8xoiPqgiTve8r96ZEnZHcE5OOL
btzSXsBuwMvsyz5sIXZtLIgLdNcoGBUNEgdknzqM2iyBcGbhD+8sNOign+EpM88CFdZ4Od4xfyhI
rSMeX5peXRiTP2myAWbiSFcumyI/9Xw9D+W8iT95MfH0qQbBea2jYuL6gWIEdvu87+vei+gxwtNs
/BV4KzRPg884w83QMw1sOyPPavQ08O5DLRm+wxSAvlC9AVAsiuQPF3XjoItZaN19PTN3fuI2z42m
sn2V4KKwkpo4N+T6Gz0JCyotjwCYllGeL1u3579HqFs/xdwhrw3zGWNexfs3UIzmqu3rdsKD94Js
BBqAnNtycFU0rhAs4bhgr5yzapArb/KokI2YLBDLxVMukaiYQiWR8FinVUolIFSOB3/13c5Oyt62
EqDkjJ+/AYVeM4b2SxnqKXOWBOM3Sz7oG0pB0rxKRRTlq3oKaS0Pt2FucWveQd6Kl3L/bW9usFSs
0t1WDHjSjAYqPYNSyYxdHvtV0wj21ptbS0a3YFjmYv5KWvbbjJjWnTB2CnLduSqc5Ml43juDfeGO
E9yz7LANbTiq8TK1hvb86WN0m5c5AOyVSVpJckl3RqlfOq79F6MrgX2MjYPF2avCfiKOyouFPIPQ
286pzSElFbEIjaDFPt0vUOgDoDOTfaKTkKQOc5lBhK/J4YVI7va4aEt2Qp6FzVuqNsYLc/0dwg5q
1T+xVLI6KJkF8mnfSM628qumcgAq7Cb3GpMlDNgGKK5KEPUNX/xhHEtHH/8JuCDc9HydWGPm7/yy
TnBuXjZJcUcUKgeqkWNNSWZZqueHFI7/3htGB0IFbWLgZISJWcrSuBG8FdQlberEZ3fxg3kk6Dy9
GqfLp+WQLxvQ7z2uNYJHxpXnQDnhp4gDlkqQxptMIVj4NJHh5tHVzT1HV1frBOa4THdkmHRlvOKl
tJaol17QIy9clnyy85gFbrf2ovwlZNuFeQLccfucDRhkfHbQ8mAGjikMtoREXnIbriXNWF13P49M
Xl5YLHxuNgUyYbN23dptlDF07Ipwrg2oJUOg8gKRWHBylH1AKO4D7DYsI8JCRKtcXJdtjCja4Lpi
Q1AZwWOSXKGpfP9bvazmHyYaNTyQTWdLUBe5heIqbG5f74t/Ctxme1O74ASrXNvo5BOuvOZiNCuU
2/yJgd2Hsnd1RoKCELbuuL0TJiVObnH4X4sZou1IEYx2M5UiFumGN8/bNuvBzUzn0SMn1EHSzIvO
9m1Ecq8fkVERm+7wDR5LuM82ARXVTQBQ1j+jV7FT7Gd2eEggTO7IcRI2exfI/YZMkDp1DBD8MEmS
jHJl2xKdHfu6ZRm2GRUWZ9xrLP8HtndghUNSN8PB9EeF9wogCPnvTaZC1kojFxc9+1AIVIxMi+bm
g5lbxREUBRqFf6om3hfMx5v+vEC8CX8EqkprmV7cPlmbYEQJJ5AqpA4CVyqtu/dZ6+hzZwhRfN3q
p51vibWVlNPPlzAh1DodiDvHIOZ+sT+D0UM3iMSH0wGemyzZ+gSilO5cHf9Zyt9s9L1Th9pemiH9
e4SrxxLpWEpccWE6FnpMv1jQfNj5RakUH+VJNTZ1AftqdaRote1SjQgWW2ioU14l0HTD7bs6E7+y
pX0/sgvDO/wYYuBs5SWLyTjaE70w+fATsbbnGW6Ry2FnKOypoGD4jYltyrbUVpLKvUf8GPjowQhW
XKO7zsOBpwoLgNTGargsa1SEt1+1rHhLWQ+svstwz+aMBL/FyPh44Myrw4pmavybEZgtykGR4+x0
sNsw6ukm0j1QIk6cIgoAWWjalL/CpEW8P4mLcN3CMSgCEdcAD6ksKqtAQ1riCB0DSpA0nHDXsvua
lFOHiM2JZX0alLn/WOXtDrJTiZOGB7aoRKIfdXgvIze6FsRWH/emlAkkuuJAzlxqtVGx9YkXk2Hr
rVZLjy1NvN8Eb1ygI9eB0q9/Pf+LXYC6ffv1DkGEu11lk9QXWZUhNsUiMuRX/N2QNXHJfbVeMiLN
qbXWmSGK0mtj06uEnVRhTFrb3z90wtVZGU5T1Tt1CssfB4bn4Q8pK8Y1b0+uKW6ixR7UYgJXBKOn
femxWVfVyWH5zlE2F9TM42BixUq8i35s2gfRa7bHBmptb9/G1mXMRuEz86z9KvA7GcId7XGcMcr9
KSwAI4LR5eJjZohqutIhqrLZwUZDrwT2IV2v4CArFPHXGK3Q/b5IfAgrIxGl/FWsvNyfByAks/3R
w9WxRmB+EAQsRlcS2aJaGpfCOJ94uJmP89Gl6Pxcz5JChLmV12pae7njNEsNAQ2kwe0TKoYc/YQf
HeoucMNNCBWG2l3XChqO3rgL6/LLPoFBivdyPOmkVSfnIQ+j9rf7NU3nizRfjxb92lyve8tvhgdu
6DdOw9XTAF2YoCDZnLHr3jJCrkz+I0LBzh4vBrQZl/9AOs2B+EpBkRJ6gBgz0S/AMnU1V+1EzzQB
CcMtXbwRozrrCSP0h6beeRjYS7Ab91gfOKbL/HiTNEhjUUh1TYm9pvFC6Yx2dxZ9s5ebCXwI3q5u
qGPP8AYEk4T5IWvtfdnI2t1QcdU6nnReSaMKM5KNKVtUC83W/J6toqpRzlX8t3DQLyYBZrMf/WfI
ssQwn2DIukW9eMQvof57Y5ID+2wP4OjyQ66+wBqIZlM+gT+TOALtc5xD8DsawZ9R+b7pCDmGGNr0
FjKYEUlf+KF6oTkDuA9dWND0csYZqJqmCc72qnu9/CutT/YiaVwgskGLRYBekX7XSQF0sbeWZeJj
TKxkIibqhl9V/m51cTFfG7QU1Mnz6YIlWyvTGb90pa0nYoVXqjw+Ck2HX/00JkEY14oAlPYnTanL
/cZAAALOtGr0uWvZ8iUuR7jk8C0X9lhS1X4J2VGhsZmxBtuBT84qi4QqsYEn86shGm69FVA229i8
ig0xIFGfi41lyboMA8gRAqwMdVyw1K/YefEGD9NaOrOSikh1G7IOCFg3XT3K2Pd37SNqaepITOP9
DDo1TNm+Rx/xSf4R9BDbw8pt9PcHagA7t0wBngMz0LymtzBqSS7l8AwzzaGYg0cGM5rjax/6luoS
B2rAN3Z29Rg4bOW1fiMU3g6StWZrDlJMqtlsQAUSNT5SOyMZe7h42ipxTsadkKnKySxopg/tjQ6o
0ONLzeqlLjpyrndMbLdrePKYPQiuDqYj8ZimBQoRMMqevTSS3gbRx4pFHlV7E4GCQYY2KD0xh4w8
CiVOOm+67YGiZJNDVL6QzXOGYqTyBxR+E0J06IWQH3q7q8p/aUvtMLjTm4rFM+di5VUjycM6T2A6
W1rk/4cf2BGUhWm/n40gWJxbEdrxzBGevbLL0GLLq+W9NcZ9Bon1QEMOxxVtTFwjGv8rIKNzQs2V
XaF/9iVrwEB3v5Eflhn/poejVSa3nRA3AklIVRGlOIjqYmQbIBXAB0NahTEXPmuLY0j1ubkcrnAG
3H9+NcfRC6mFXdhKVZCwnZBrQ2yekeTO7CdUWhjgz0t5mHA4SWhwdHe0YEBs2ixVikLqixuoYK3E
BrE/z/B7uT7NbxHB3hKxq1E1jPc3z6uYqpys1jRGZCMqTgajZX/4D1CWww7CNf3mzQ7yc8hNw2Uz
BL33FTZ3CO9pqzgMMp/LkhkzysXlNjrlqZHk4DRmH08hi5i1J19Fh1SkuwdyN9SP+AWI8ye4JORy
9RQUwe+9TXQ4GU6EED/t1mNjgy7LUA91qEh2+PkPuPAn/uY+QfuUnmeJBa+LiuEZ3EkLpba172wP
h4ZqXMdW/ALm2wwbuqqYgH4mbFsp5SijaogjbDhXoGeVJ1t00wkgHzzC8R2CKQjzsQuRbW4ko4BY
bz4bcLgo/Ve1ltxqamyZsfgwlFlkOacrBDvOvQDNdlIT8ysggAEKXMSeqbeSkqY9URS5PH0pilvV
dgsA2n/wTGjgbbw+rTTnkDaMkIfLqEU0QeZxwMbp8ZwKqpw8Rx2m0Rkio70bilLoCZy9c/YJ7jPu
UWYKBF497VJarIoYS7tykqiPdrHCWk9EqV111rgY+J8VnEieUzo5N8Cco1NbdtENdvesvRobfmKg
bOXmj3JWXGBUdmatT9zC6uJbeLMIf9cVCEOIN+4sNW0DTiSaX5WwiSujlvJBIV3fMdWVj9lb+d7s
NRpBSm+Py1FGG987smEwBlzIbdBQKPslVs/Dge2YJYwJrKLJbIudUfQvY7uMfeep5AvxSyDellIM
RrvO+etyQ2ikJGg5uRfc83cAgALSLAWqe6lQrhZ6vQNoeWKYkaJdI8RR5hAH+qW5nYb8u9e1qz4w
DXvZBi0GT7ZyWDzW7hV29hwSG5nyLg8KoWxgDcdl4qhtRnEaC0HFgiW9hW/K4G08umB0b9sinLcI
+NNz+0/ixnkHUf4GJHDB4JtjFldCfHiJJs4l5sIcxZTYRsIAq7q/sFi/FzIxXTUxZ1hULazBidXp
ZvKDOR06k694BjMcJR7k1hcUNN9rYUp3M3/XuukAn+Y2iNRnDMnXH8WcTPRIhdvRay6/tr1E2vub
uOPC0UGKRfO5929SY+nVx/Z2WQ0pFKuHkDCdQO+a2WLpz30VBVj4h94h3yXTaZmQsZBcPdzqvDbD
4tFUYMcOFT+xf0WRvXtWEgu/B7VKzNZZWaRfNTbAd3wRpseOZBh3lJzHLTE0B5V8lnzt3r0K/fHj
xY4of3tmp9Gvd2/SdubaVTQpb8PkjGJrRavSLGArMWnJ2gujtR3YglCKo/5gjA/1RTljiHXk4NyJ
Syd8NhsEE8Aamz0FuY9GXhoX93ULxwHe9mFYxy7nycaWU+jxlNeKXfqOSFL8xUw9a7ZgQNMzr+2Y
+llPAEqvYqYG6MZ3Q4eZIxcK1VWHl9/79QQXh3x1m4bMLikvG7eOcs520RCXC2sHM9OSSGT3rDTj
9XTBNVDjGG/KYFSOoPp7r7ruLopYSbL8iQXYO+bjN1K5VSDKtkgfPDEJp4/UFoMGEUelJOFGo//G
n3S/RadW/yI4LY8KfJcDlYf4RBTcAsIddTihhAA5Ga+wQYGXGWt+jSoBgHAZJG6fSmcQy2ViaP/r
fY9Zeev6fRhLiTFxqtNxnLCbIs1LIHQaErMi7OCQrCMrJktak5P/TKF/Kah/YtyRwnFBsqcECaPB
698sXJJQlKPsG4rLQgh+3Xa9Q38jmkky0HSrAQi1SAWSM0XlmiaKwfo0r769Vq8Ev7E8KrzWOmwV
EzhE9YjIOQAlNZ90FEslBDpJVH6Ffw6hprKdsG3nhNbeBp6chOiTo48uFe9f6sGd+EWocCLOP4TJ
bYOE9eu6nnzWCfp7aKj4bH+IFae5yh5pnTnkPsghJ2LI2RsBc8rJgbBXA184UnWQ18hBlV0hk564
pWm/HJV+l2IoHtRZYn/21IGnWpVYNeHhOnbIgVhklS2Hs1xEKGX9uzy3EjdT30f+Au8P9ryCtJzP
RVSg942p0WpaXSr7RIdboq/7IHV0Dq4vwpkOJ40XKohjTQQZEYNjkdBJK93+nW8+GJNjVjQlvF72
JjVN/FID6lmMKK2Xmq+2tbiUfu1xunE/IvAJK8FxMAthe3iPYKlXDTiyrdw0opq56XzE5kQutBAD
ibBl6mGvnLi0ruje5IMR0FOHEIlTd/Y9HRObc9vRItJgJdlbhwSh4kiFmMceCpijyCUyEIivuxoR
FcIOafA39dxyzG8UVk7j1wMnY0umdiAWwMwrW5aE0dOm/WO6O9oyXGzPNGYxazZOwdYtY+hZH4hJ
SBocgfbp5FYrCXD11UXbZJfiWZ4ejnCS03azhlGAz6rF2Wj1EKbjZcUB4SEXG7pCercuGdFM8LZC
cFlD0BZvX3DAJOsnBkWQhCuRUOtYr6M2XXdqk1+3oFaBoUm+T8akn8MijLMMCQ1yMoFkGR2F8Oqn
xnNbtd4xW4Qu81weM0H2YthCsyt1opEDMCudXaLk1PzFZhmtIZTTUXtpEB+CbE+5poyhieQ2cGdx
K5Fm57FGYY000rqjcYoK0ZZVuIbNM4/j4Zx7eNYFCw4AjF6EHxpgds1sdxSy0N9EXro9CMAlb9yx
zVAl+onZXbthmG4py43Si7wGtm4otXyhN57dFaDJNOY2Pr1Y4eKmNaimXOZgYEVybAanLO6vwUaw
Tu1C0ayfLxVDb3MLfiZPzktjViIofAYsEIiKYyuER/dQjQJ/5kRFpYC/YKM5QzGeOs+xPrSmX+21
4wIkxcfVpyI7WJDA+OzJRtggCilRTGGPUYox2xKWl7TKqwK/6N5FT158B5fxtS4Thw4Alk72fs5R
PoeFcz+TqJDhBJ78EnrTE2fbPuor56rVT80g8uA3XtEELaASzL0vVf75/k4re68wXCiFXfBPY6PA
BQtNlt1WAOPo9A8Nm6gz3AE203VcQb348gx8WxM3kS+44c/EMyMspXPLViMpP41AFRB68CuZjSxP
8ma84BLUOyoScNB9P1cyEudSZSmC7hTTkC8Zat+oooNbQdC3tuwQHt0DL8yYs+eJ8pXgFpCgu0K7
DJzJDpl1+uSBe/+ww+R57IVHm1S/bSVN2EPlGomDWKCr1otXqd8yVmjwfmlDQKBJmgHtQnz5Gfxb
FTLLCXizDVw+ZbO0/KDm2pdPpjN6nvhr3KPPHqpnruTuM0YPNV7fHk0c+xiDVEjhPsKvLttkHhjG
0sSMX1kh9Y1h+pLbzglqS2O0vBlbSOLgyxwSACTKmf5ngjIEXlAUfGrSmxD8cQPhmvfXpKgenD3J
uCU8wtJ8CdMYxtnqGJlchWzSoh440JB4SMakAE28q3FhAZMiCpprJDL9U04tDYvhnuhEcLEWe0vS
vdvguE/bXIRGv46MDTiF1MajhknTvCj1bKv8Kz0nOMtMX0PWdUUpQCvmnj0fZTR+w9NkFYsNE02y
CqdpM1sR4klWDwTY4pTe9ls63swgFwTGKnGnwyy8gAsUq2aCfxrj/pDK6dQ4S+b+qnq/eeE7Jg/n
4FD6IZzHaIZchYllzT4Qm77BeMib8Z16RlNZkPf9izHvSPq4Vi/PtgHgF6VKA0P8sofGdWxq0onr
jXdHRdSWDrTcEykL+lQ2t3E6lC2YC7CjpbkFgSeHBya1pgrekuKYgk9hihB1ErawXkT8VdT5OEIu
vI+6N9sW+H4kkBhWsT77AgJfEz2iilvNGg3xcj/JuHEPxsAJLYeWM+5hnU4q5JyeMJteQBO9qfAk
P0Li+WdLfbSILYAIcAGFamBF61geMLW95d19y0GWNoERPOPNW95f5hpM76n/VNIyB4dc0WycwzwE
nCIQmmtXByB7YXi/3qQNvB6lofBkDTrm60DaqTDVP8upe7npvEbkFS0OGHh23GQJl/Mn+qnAJqnJ
sjHKLuIAEi2q9dBjn+0LE/8uYWLjXJ5lAta5jY+Wxv/8BSFsNwh8yu8IhzOBkxPe+HzT8aw6FSxW
qFIh7enw6Ft8I+ZX0zfbGa2RRkqC8niRKn4gYcmtALowkAjTxQz0Wk/4Zk1hC5xbkUKrzDZrz9eC
QoBt3Vc47O0iubera6mLTBHtNGxOn9dLnePidqRYYYJnonHt7HHKgiBu7fC914w28mBUxh0DTyT4
xACjE2qmN5UDwNOZEIn9g/hKznh7Vqr4si5wP9TZsqQ4lNt89EkUURfQugiJH5vrw0dUltkxtHKe
F+CQIXB8D081/7EcaroNXIUXaFYOepJD+cKWWF0R7CRVcSkFG+U7WFEvTkQ1XZ1yC5jbSfdv7Gbi
XigYVe5lGMkDMdxIqE9oFyR2H8LkeJBKTnvdTLjABmLENNKU2ASzDvF10xGNzmoDbr4Ez6kpW8rn
KC+5Yaza6aunDGsgY6G4l7+qiztHx2wAA5l5PiuyaJB3yCumZit76/rNDwtv9mdYDB6FFtI0DxnM
ZNo8jCY6mYEWAhxWZI47JdLaLoJZ15qZSpGpSSs5KyOpV9EeqDyNitIomzlKesQTWMT1M1NE+P91
oruQ8MamqZuMeryCYNaWR13HkgF+V9hBu1srgW6o3Q+RBmjGy7Ju8ncxcuslOc3odvcA/sfINbxg
VAeMXcJuYdN/nX12cpM9XxENoHp14p3VOQNdQeCArR0y1dWce8UgUkJ7/b2fUjE3yGTaJHR6WC6N
TRLv0fCcOF1Ss8hYngJStTtvbFo2S7Yq+XpvYF4Qx3cnzSRwFHcMkftJOO6O/jSzxgsoJZmnLSvY
7ZNwfCaI+2OVUQWC2rMqbSX8o1XOmnCgdu5EZe8xrVm+GxkZrqZAKJiuukqi1/IoUUQjthUH3b52
39eB1gkjIoaUhay3an8vzUmMTTxSjumIV0Byj14DUNPxSYkxJ5v4nRg7JwJN86ek9oNKA03I3ziw
aW76Wbu3XrudvHYSZS1t8uzFXj7t+EcS6PvLH63QMarrIbkc3aUhMvB/4wyoA7YLeXlEKzHPnxY7
5QQdS8TZh0Z4+nh440FklHNQPoxN+LCDtUrY3NsQTE529kiSkpuc+j5hNuXyaiHjX160HYZGrTMX
FF2Sv4Cme08eBk3hjU0kUwKNOVMaZrpOGE8tVF1OOo0jdPDz/oznG/yslRUBETptOCII+uGKbbCn
qFnEW+18XBEXdUo2+H2+HyUpO2JQEJfKnUIdIQ/+ffV45IWWqB+OuRER6Ntne7hlee30tTbdcdkF
FJusTfikVlhQOljBotwGjMeBdbLDjGK+xXCZTIEm/ICYXz4vrH5b8M5nys0TOzowF5RSTgffaXEH
i/F0u5UTVSKIIV9DTcfZ3gMPCuqvYuvteUNc9HXqtK9La37X/4Mg53xrinXfYqSgLHzno1H4zt0U
NvSLuTRr67JBMCkesrBgjS5VFDdQtJY1KQq0ZwB6qIG6i0NXB1OJhGbqJ0xwr+KlQ/yY8q+TkY4O
vMKVI9dnMME8rpbtrDGB6/X2peKRpPUoVqp7f6G/qqVO94+fWZ781n5YFKlm+DQ6Ok8kwbW9qpu5
mk7mSJ8UDisr19f7jm+dQBWJM1ktfyYhHCuPjYUJ9LYLReOgsQfNUsfZd9dlT6s0uU8Ip1zxHvZc
Wks8d3m+iaZuYUKc3INcRV3E0dxksPhut8U9h2CuxX1yN9XjhrVw0iUq95V+WlJWx9hFwV/mOzj/
ZpZW8eSzD8j+GVWxNKqrDeC3soHMZ5WfeEvMNJHavOcAntdGdzqtqnfyKqp9G2N3ASGuXRAvW+rK
T9p0c0zQmvz1SeCx+rlPhIWNTgW7qksRbvrJYy+k6vgaIS74r/MbMfehwYWnKYKGtn+wtlxrWrMk
wy84m1WVydhJytYsjnIlf4IHqwsGVDH749FRI4SjGb+u1X/MCgGL5Ee2ufdxOEgE/aSvSiw+4zXT
01hULsrDp96wQ/QNdSFHBjN1fygRoTn2MRmSEQEtCu0b0mio+GRHWy/sPYRsRU782VyFYoyJjzXF
k23yyM8G7ew/T5kbYr555PGbb6lYus2vlkyvINp/FYQJD7cnt1NBgUXGhiGZUnvVbiwJFB1/v79G
GjHvcYql9kQPSj73c7aJQ47yReAr8qBY2Pzl+8u+88gKV0s2B7v5kG8+IvqqSMY3opBq9wEAU+EI
a2gQ5Bkb/tr7kd9lpf16GKS2GC8m3Z5LpvJ2WXVHrJ23oMyBJDTkaVw9r0VQ+Y8zaWgwEe8PqOzJ
WqnGaiRxABH1kALS+KsC2ahpK6DLFP6w2xJFDrdcEhy4ASA8FR1jqX9XWT7xKMUTyEzWxJ0Ip1Mr
+sZoXutBIt75YcfsZKgntal5yRivEaXIex9AUOl4vRyhf5EqD89UBLiBHcDRagkcbx9ZblxJNYNy
UtWtbts36uYiP8YLynt2BDCr6ycvFnfiv1d9aaOb9+ifYX29nKQW1D6SfYPAU1i9/tBlOH9u8eek
aMUkndyHOKHaYtjgOHvo1v4SDCtEZcKSYmo21D/w8UKzk3zsxoIsAPzM9f7/0ojxgKQpkb3bHubK
3BwGadgqQRxvU3DxxaUtqg4YCl1bafgfPGGl1v76qPNowZ4qaaH0vHOI/O270tjoT7uQCiMNYL3V
DTnDcSjcakVT7o7hO1W1TuRS4L5sE045MbgD3ziVtL0RtwFKr+d7dv0ZWkTwcMibnvJjPxYOVJx9
8Lk3NF4jKs3Ld2GGUoIjEGKPgfY0N2jxvOhmdZPRREBSttOCaUnc5bTWg661UwViFzYpPrUlJ2m1
1QSq/jt7jYW7g2vsUwgGaeioxHJQ10wP1Ry63Hm6L8GAD0Q7PyvgibvdzCls62V0UIFNWD/pEsNS
Apop3LqeZAsCmD9zcu0qfpJjsfSolQIC/Hl5kHFOD3r/I5sPI0CZEncVoC3tR83Zz3Ty+Ml4nfCj
2HqEHj3jXPu/Fo5UFYwE1fAH/5y/pJI9pgGKXRtXXJXprULwxLsQW4q+f3sStvbGzendeTs01Ibl
RxuE0evGPuIMwuNzzN1lsMPCW2al0763fKC95o3daRWQEo3ggXENWFywaGsLE1734y3Y+xL3d6uq
VI4zHPpeJTUj8zrr3PtjGSl261O4+8gf9vswMb2XZxEcQLZrkFg2hs3Vh7dH6+b/8MiM3o4DKhxR
Rs/CAXKRJOLv45HM9H/PTRQlvfe76UNpHmyq2+Lx99tyUMfaSdXUgTpc5Sfwcosu5coYHpHIK8Sy
45rBapBTITQvY23G48ni+WvzVbY7DdRCKVh7O7p4eu+VBZ+MTn/a454m1j/vhHmqnIUq5j1WodR3
VlUvpCLg/doV1eBMqwUSP+GoAqxd/JbrQ3B3jux40vjIntz7aV4mbEgnCmFg8Z1zXoD1W1LuTYBl
/wUBlMf3/z0xBxmX26sY6hkMrzjATpRXGFk8Z4torCpYYWNPpz87bpbag1WWculwxPRODrG6uP6x
3Z+N5yGY9V0HjEYm7cjgF7Rhc22n0AqKbrkKyMZpmhzuSztgXwPhlDh2jWnKWYLX38uYuPRS8p2/
Kp802+MGiNOUhGKiBOyAEL2BQC9q0hvh5KmII9qR09vh/GkQiO9jVOvtf6TCQ6Jgt1Kyc4VGmm/w
RS0JE30kd79DeRPgHrIFD2gdre56GhIltC+P/ZNrRrYh8Jd8u/I2jxA5Ej8dUQpnEdy6qSlHubCM
ofJYMnjayHfjo67vzfs61/A5owPeGe+AhPgF7ss9107XjYragIveySsTRYgID+Il2sm23PJVsNeR
fKJcUoGnPw+3Ny2o/CYXskKikv1UzNKDKiD8hffvgvCk2ugWagrmYe9V47FfvLnq7uACHs5+sCFF
9Z8gDL1LJj/Y2mFWvAhQQFZfjlh+YJlxY5HdqVUId7UG6zgB7DSVOFwpQ9KRGFdC9ua6/C9ewTxY
1TsvstA58Xbkgh0BGbmue2XhIm2Ck19WWDU3pgXRYcDg9dRiuDVA0LEzkfwxG0fx/qrqCiu13qPm
0s+qBHbfhd/ckXIpDkJ+8hfOwV4utyyla/Qobpq/6qjKdAvLE+FKGn/yoLgL3jVVnnpcpADc7Fn/
Y8IQh5ZeZwlPbB43ECVk0VR/JQ8ctXumIl+3PAt+u00tHXw77ziMPS7+Lo844co0fyjlzczjqJe0
JFb1IYt/+3mcK9oUj2daQE7lWBHekGYoA2wEGwHvm+9rfAfDUcnT/vFybg6qraHTngRfQo2xvIrM
SxOi4EfrkRr4eXEfmXLXF83fm2iNATBgakntzDEpt7j9do6O57o5TqwAH9+TCnvv77TyFp+IRTLL
QqKJvffUcUw7H/DhauPe5P6xXTJGADLKd4XyXrT4EGkG9cJe645nUIVRuwWgfGi0FaPfZV/G4hlS
sbMVFsJwfrSHp95Wdqtxf/YRxlExhQ/XpFhT1aqZwWb3sC+kKRIfeNjoht0N2angZyhnI5/vSR5C
HPtqxBtdzFXIoBVLWdvTDnzK2zWqKuX1iyua0VTWDYLy5lSqX1pAdP08oKu8KI91xBDr/HlbBk3U
Z/Bdizf9ex7bzF+QZcWydvva9et6fvVBVwfqQzRNCCRloNpyaT/eEKHa7vjmLXa6bQBX2/B5Ql0R
Jb64rRFxUU3pBgvQhJYCSK2+JUnppn4ec9IGwzf7CLvRTjXUyGhKDxda4Jt136WVhgwgr85xWUdK
wYAhVLftJyfKoy5fVzZ7HXNdGfzMJsL2P9rQ7tP4WUc6/dKh9m7viWawGmriX0o/LZDm9uXvglv4
50kJCJ/nw94XyTaCkw0FyC74V96csFCV/1fpIHkUAIWUXBtwzkgVtNGiDSWAyF/WpzjtGkGt8Rd6
cQ9ngA6ashJIRaXI8aEkeA3AbhOAIxEFZoxdHy+yFuLNbE4piLVYI8axqQ34H4Jz8ALOo8jIJVPY
ACw+nY+EJxx9ae/W18PZVCz4i8oLaYN4o3hzRVEJgCg1ecR/NZq6ToSFCVJSYpXmDMn+yG2+BKO3
L6uigdKKx/kLlqHKxHYfPaIoGTWY5AMn7oXaEsZwgC5y7DMyh9mZ0/W0QHHPtR6KMaZUMv9IoJ/s
A0yYxD7objATYg16phqXG13Jpo/A4r/YvErCsKSKfKyW0W1mHnpV2SEADrZX7JD766X2jC7CKGhA
Zw3O9oYG9/lbGdaI8FUDPZTisdZ1mPfei+34Te1R6bicbF0xCaOGwLQcMqeyjdS92JUT/9mKgeQt
Y4ooora9KskKmKK6+OhIMrZ4hqm4juz5dEp7vf71p44OkAVvEcO0giOPLIJ3T47zpk+lZ+b5XiWZ
KyNaS4sTG9dJlJSbtiEThVDeBtMEWPJvFMGtVPrYC2+X6SRsf1k54xilnJKqc0MSdmCQnK2Zu8Ek
RtBx93h7N32f7pZoktB0oCxZHIT2HBYfOkvzK58mwOPDXKSXNAUy7a0awqM5e2H2bbVGWto+ji7l
ncHXjQnJ1mUMcKNDMchMdK+4MABbDuLHtDi0wwIr9g8AU5bbt87RSUi8jMYUOOcbo8XtpbgY3cNp
3JooAeAIggUB26LkQA3ngk3h5DQuc/MDlSUONO6+PQp5zKo+xxByChHqb9R+RaqqIWPeArga2uH+
iHgYrEYePemcxDewJ6prlA+6sfKos+MI3zMW0GkLlPwxV7ELA+aySb4dgYLZQJY5lyHyrwjNNpGE
SVGWAcQTmiSsCq1RWlw1bhl4Os+UMbzCZAiZq0gyP24Mqs6DojfyI4Qfhr7OhT0Azd3eWPXfMY8+
0mHY3yxr8Uh77Wj+UYOz0Cs93+x16I8eMp3jnbU78dFF/b1g67N+FOwZD+7LJqTsVp+1LS/RRKeP
jqbD5DJhM1wNQO40cluV6eOgsHiIATUdW0wHKIvzjmOY84WIEN7UdZbxbkOSCnWdN8Gzq2ZGD2ZB
XTCb24SSG4ziSd+QQc/FNYejWEicVjwnfS4jonsD6N2r8imiUliysGauVR6vNRgfZiywIMNhL6WE
c2ZgM2iWr2leosk6PCLtfXVxbt8/zaC+RNKt0iUvJimWyzGf7MFSOboyHepBdPzFnqlRwvI66KZv
lKBmutiw+3YYKnNxTiVHi+WAFV9u80c9dc73DVsvd/OufwffyVK6slw6Lb+Zs5+gABAs2apRbEiJ
UY7ZTdSqBrjc0jRjTMhJDfmJDTjNaaLhFIwKiFFy8k2NF/stU0O1aT9WIx8ZGqjhbZV4Lia14ju0
ZWP3rEhdIfj9SNlcaE0pw5kj5c+WvrThEAUZBaHDvNuJruuX4uCedksz5Og09XN71wTLn+OtpE3k
k7mfunJ+Ar8FvEEZVSHBQUQ+m5JwH7BIDs39Hri9fHIeW4aMW6dWsU4KC4dOs/n/LnMaKtvNDzaV
58wOzz7b3XzKk9x+30dXcRp95dJyvzu2tH7LejvBhqouwZVzWzgwazP1svtVhJObO5Ff8uJdJW+N
v08X9/ZvHCvJP79zPfN3HuuFEBuq3d6hHP3WxmTjRH3tUJ1wUIQUMaD2UcaWMn/Gnu58GDaTkQUT
Vprb5P0fIn7zkqtNNoB7vO59XIe1t5Lp36VavtlrSC6JrRoUQzY1rLmGbk5EJJsk9Bat3gzNuloW
zdM9jDK/6MYl6vdJv7fkTAdszGfTI0XZ5XtH7vGbxAPtEIr7OrIgMEX1HJJqdPa39EcJDHIRtvGs
B+dJKmcsw149dVD04qTvGPrQ9y2utA9S0Hib6rYmiW127tMW/cVdzzS9DC3PLf6hL5DUp7HTwmSa
DPQAxm6iKYlxrGH2K6FC1MEWqqJfCi259K4jq01SAbOlIPB8ecz9DAKwO5xgr+3fgMeO7XgaRMAc
ilPrBgDoifYA1ztxIZaaSprdcXuxmsZ06F7oJ+ciGJgauSj2l7I6SAYH6UIsK2xSTVQu0J0cXBff
oag6mbZSIbLbFfDCMP2/ViwWq69LYseOnqUta5PlqlTpv9Y+lZlz+vFZcYnesxUy24vcM8xxhMhE
H6n5wE2UbOf51MKNNRgXqaNL3InahDGiVJcRn9jyuq5HW0KnGoRl2uBu4Uh1wJ8OabV3C158MZoG
/aMlCoj847N4ot2hX9sHlaCHAyBugxGfJbj9DDDhWeaJ1yxnwcH2C8PmJsmH0Gzk2jlFkNwU0nmP
/IzXP64q3/Ee+bkJ7wlRhzP37vZpOa4O9CN6CNCkiqP99auo5ljGFAULX/t6lGi7aBg+Zi6f2il5
iWckstU6YEL88oOB01iZDwkVjvUhCel8e/8NO7jjiIdtDslB+bwNW3SNGwQ8eJ80SbLM6oQeCsjv
cZ+8mVfF67EGYjEnBDo3MlEh06Hce6MM22wq3A85cu75dsjzjLZnGfsc3xv6K/dyncmui4XXlPpH
YPQtgklLpegiPbQYge7ZwGUV6hnSkQR1jgdPGZVT2v2vDh76ZNt7DrLtsDbDXKFRSm8c/VgHjJrA
ld3ZVO31ttp1LrZgMIww/13GiNrX4CYZrVC0EhX6qX3EiIqP7H0GV47vR4LEAbjBrTiVm4vCyKji
jePHR4fYS9g6GBfgVyQrADnVMawYGKbCOdjnR350c3Fu0GcQd4/47FGFWk1hcDVXYpyPwt4m47Fu
uG+qlzE4Ol33tYdfM7fRc1PlTgaYIT3sO5AdNc2VcVqeaSY+qzf1J+vS6giWOKfEkhWJp5SZehVG
fjk/iV2Xsdc0owL7oBR0c+JY3tPvFakT8//nEkoAnD7L7rClEYc2vLJgT0cFj4kp8cPcg/FdNzP3
fncSDkfWmHzKu7/zvJSqgtztaSo+oh55tYU+0lbQgmFktPxRgZur0KMDbRYOL0RF0G7kw+qypYzM
pNWg893hiQxhENkf1jZWDoxRmdGxPqTgnZiz8wNtCP/IK9D/et8LwOKJcF2ZC+KXjcx9dd2Ye9r9
QGE972jVrlhzQGlr21uINt1cI5gpHy0QKKFZrPm192jFHoS1tdVLphOo8ouNx62bVvnQHpGr76LR
rfMDlVQvQqO/Ehhhvqzc+sP9NJDrMIE3yUwGXHDhSbnCWzi9PglM/B3VSdjPRBU8SbYYBy7rBdOn
ZRyDjfrLq4A2c0oS4pNgZzm6UYQqEXx40RBvZ7aaFG9h1UTKK9mOLmJI8kLP4V35FmfAVv7i2tz3
T2wVmvhk9q0hzc0eAGl25+osZAhyg/Hpyv2yrL4eN7Izhl5JxtF1mk+GEHbx0MCWyH7iufydDPgw
YSxyJzchIPA43CaKWvoOFt9JY69azpnNuI88hIeBWBLyzLvHlWlRdstLRRw5gRGfGsD5yvfV6GvP
gFqOpMJDznfXXuTsuyoZH+8mXlnhXdm75r1tmP31f4L4Hz6Nxx90DyG106tFhxrn+M378kCpTuDj
rXD5ebsJKzxe1F8zIhbNZ1DX49rs2StpviPWzeddb2DpFuL0OJnRdmO+uYYeUBPGXsAXYUhN+O+0
BQjegZwrL4dmuqFL0lLduDwvR/2UEJVREPYAzoCFmPutqpgnORGNBJBlag2wivYLZfMbKol4ehU3
3WwMw2n05hALYWm94ZEB4i1rZ38doRAtsfedhCS1F5u/L2cGu5Va/6GGsxo1/OBXYNB9F1UZVf5q
GtLqg7IWJqq022yM6uESuhaRlHtEHt0abOpV0cOHR+kQUenEwMewN3SABa46XbtRZHDxZyFR9idd
z+6ii+QQ+68wDY6JF21peUvktcuv3GhLqz9+SIEvKS+HfAKlPsysYAtNfgEV636NheWnSYa3JHiV
fLkouAC48OI0jrqgI3CWtzfK9IHOqiBHPE4ytQ+7qKwJ0w7oW6vM5jTsB9BbzEf7OtsZmGVzoy83
rth8prCeGxxRuNvYGehik+rlJ9QMjhYtOyPqSZhjyPt4HWflr5Lbt61JBbR2XeuDjhjP59cxgHEl
GAWnOiC216g54xXEe3k42Z1eFevuLdm6pRK5kCpkQ/UnYdS37Dt/24oGYQ9eXpWCnXZVMGjdfTIu
F/zQNBinsK0go56ptqAqLL7ieKA+7MLyCVlj+0g1UIR9vQuJOVtbYnWEfiI5NVGvUIMyTKFVHPrV
wyGFt4bmI01Cpr5CX5Y3ObiAR2U1BAbmrLhRVdobJXUOpz0JmXd/k7elsJl8c9xr4qDJV9CtPuy1
YS9A6d3GD4N6hr2ID5kKr0tYh2TpqDTExRdRywd9dD99iPCXsEcz3OC6TV/Ea2AfLb8B45yJTSje
K2cY5RgFZIf9J6ltaERex0hJ+pBfqR28u1+oIP9s+khPpNaratuIl6BqdPce9qAY49fkseOhiSCP
gnj4f5qw0pyn3ti5AnXukR6fzXfk1MgzZIBEOayoW0qF2LnENGrvWjiuFchx78xa6WwUUymjx0Kb
RoHX0X70xd8i0br/aVBS8z4gtzdBmZyO7I2p5lKMrLJq3P7OQDUPg4CdvAylmg5qYXxXdJ+64etR
U//mDwbhsfv+Ycc7id+USGwl22YvYEd0LwrgJ0bTFx2giZ39swTP2MmJJTsG3cpG9FF5mVUJAnqX
1EbjmLcIGywF7rVDp9RP24nawtACpqn7Bn6nh2pzZ9bcFWj4+qJUYxGJWLX5zKL4/4t+LQ8eYxBd
A2yoAYb/MkN7afFYCPe1sFH3ypreOxbTYVoYrmLNkK/izw9KtaOr+PD/k4boxovTsSF7vP4q3KEn
ERsqQTspm+LgyrzSzRik2KTBfBJEkHXWNWpvCJqCg2J06IRufbBo6vNGbi84VaMu1NCXPf7k87QN
NwZfrDc9gbbgvisvQYeOS55aoRc1XF5U5VP1hD/+oXxZKg47xNBqaKSMmsmeS4FJfj+uTff65Fym
NpEkd081lU3UsG43oZfbywG/cqis1j0LJuZ2X9p4OeANwGCdcmBIbyGpKOCTxsqk8+/qdVa2hmla
J9lvDdNISZ+xYxp1rqZSreHStfKPR3+pYtuE55Wkqg1xAlR0aVzFvTVYqnxvf7j2bDPrC6zd8Qp5
FXftmK261KJmsTMkPMsuR0tH1ikHzjfzghu/XiPEwRx0W170E4BD5+8U5xujbP6reCMQCSOjUyQj
GXiGnff11h/jyb0BlZpN6L3aP8qWCdxus0HtihFYSsft9Jk0lmvQ8o1OuqKRiF5E99m69q+CqlPE
KAv3yECpb4fYhXjdfKPQ1D1a9+ZVW6bJdKTtadzSWQKbGBqhz8c0hJM7CYGs/YZAsd/diummXKYJ
XnOSoLJTApKcN/pZ1Xr0xUzAJ5yjdW9xy+QFWa9AbaBhNRqTQ7CYrTe1z5LF2Xfqwoow6+cPu+FY
5fuqdmd0y10fX8Y2CMegdQoxNVtvPE6SYaiGmFjHuLB4AulXsudvpjsLpXWEDLfwiSUqveD88hC/
gw9F8TacMw4/ZFltVBFCdXuctNkaOlW7RKsh3Ob9woNhTk1IQlGAV3z2N7JuVcRnQ932eM+O8Ynf
tkvtN8bVE2xG+tbSaIncjYrxMLGYZELVXqUareEnQk/mTDr6LQzE0xziGse9u3NBWd1GLy/Ck+AI
sNjp6QFeEcIX/ixej88isb/u2p/4p9vDMfKyCSUgU8S+hnmYNdber28C0anph0wi0gFECy9OGCjl
aM7oixjVlGnk1jnHym0cG6lAuuSo8Qqx8oyWPzZuFzsN2fwIZ4UU/ZWS4QDLYjYUGO+s1EbLJmyw
i8KY7WXPPGlfciujbNU1u2AWPlmRFyN7jLVxzTM+YRMavtNEbdajCu26iUFmYvTTuSWfnTc/9OZ8
OHqU/b6C9RdeRG2cZffRLZo4FfbFIMeK6dAKZZ8GybupbIfso6HtHoPvRVFPlNyQSUhNRVhhajwK
TMk+UBaODMUgbsliyiriIAoXK9UinQ48d/iitO9BhfcJOJ59lfm+2pT/vIXFBT1lqa+dxPsnUi63
rFZ2GkSWfCvBgJrXZl+KguYl3VRyTcong2xXQF3skwDV9PZVp8ZoAlWIx99NnU4xX5pSVoJM9LDH
yJAAHrL97UI0FkKXbmhn1qmzmL7k/1Er/r3q+22iX82gD2WaK00FrTzRT6nwbEx7kRlBpb3AIGKE
6pvAR9FaNgpsAHWcxY1Asc3084Q6BHbwMoizP73lBj1zWutdAF7ycRfgsZPcHNDnYXN42XGN8klP
3BzWbcxa4Kv3cSwRiMtVFu38tFQYCVPpsEwEwypyk/YkyQvqmJHHoz0KNQIKD+j3vUQQ6kEn0spA
JPKpdx4vB6mCcTrrB3MMZ9LGayIMRfZc7h7boZ5xqhamwb5ScMo6KlsvxP+UPaFyyyTvK+MK1Cmt
gyurwgJ6IS/iNUAmkeen8Hgg9UaJmAlqxOSO6jvKVW4PPnT1SUwqg5Ce9gvAHRUKYCwvEAcA7m7S
qm+1etCo1ngkPJdsX6OGwnZsi1l6DyRAz1v+U6qk+IbRgbM8IfpoUhNMZDcnio1Pgu7FIidnXoF7
tJ8gwkM62ij+8WStb+4L9lH8gZa27xGc1NpAKT8o2bK1S4kXPwtMe9oRAfgA1x/imbQYEEAIW9Bs
ghurvr071NUKuUuehrYN+n4oE+iRTTyF1WbpMCnY64XdHnUO5ZNCPzBhkO4hwt74OV+syHVBwS6n
w8zwikBqOtSR/uZ9qlmnF2glr60BBGLjlwDCuhvcajSrPuGlJqPryzN7YHcTIHKwV9rRyk7uZF+e
63kQ37znph3lHznl8cbVMR65HiOIVLpRbtI82OfWWALqEAJ0BlmEwInnP3wgyhTjs3bq9xY1MuTT
DS9jP+j41UsSzOZxO0BzZAp12tcd6T2MY2Sl+RP0rJEC+cfS+T92aUqKBDv8G2t19jKSLjQdTa6o
FxHfxo4gc7Kmla1KQJNlwChzHHNQ+DUFAeioMKqZTmuCA0Dlfb0BS3oWvX5jQb7gBR5SIFN9E89e
xkoNc01U1EyECTGzHZbpk+TwC68ZRu2+aTBdgpz5G6uyOICf6xa6+XAde6QsIcohM9bZPmd9bA6X
U7JVnMc+J/Sa3/hIX/6UXnAn3qftD6a4720weyIAncBit8Lmc4n9zg3LPrGFIQGPqKkfpRGu7Sww
NpE1PJtfdiXuflYxcL4pwXvtJJ/zluY0u4WgCEVyKuki11gBZjRKW6DlmhHUQ5oK6dnQDvMBTZzK
Zkwe7tnxFrSZtCc6iM97v1WG8mmNHYacXcii0V03tyOINdiujDiLPza10IkcD6Web9ZYVDR4f7n2
v8yscM8nNsAbKx7tm0IdLzhzt1SC8KhDAdZ/3CWZ0zIxBFwhsW42XRKlKJCmKHU++jJxFY/yOjVU
xfxl50uwY4Lu2mnJsW7qgUxp7iTa4p3Fo3BnYXckGCa1lgja0jGmYTyesFyJnFcY+Quzz92S2ZtZ
nIcTb33mUpXbowf9d/c/KGcrIv2i3hYhlF/ImRzEeD8svy/UxKsMI52PkTKnv/ot0FBy3bg66+o7
D4icPcZY5ktBzMRk15v86U4ZYGriWHGwfw1LNjW41n4zb9kgw83yY/4xiNBGwK6XvW3ixm9kOEN0
7moIsavyq9gOVQjjXTPPzXDdXgOZe8Gbb/0sOXwZV+paSogxw3kKejMgS5SjK0SMJDUV/ySxFg4e
4PeJ1FLeuzbGp5tVNQ91nnZENjkdTldBvGiBAgss8fTPV58yakr5XLwV9uMUrinEMwJHL1D8yuPP
+ktM/EduxlrEbbHqw1gverlRVLMVSpxrUtKu7/HU0KzQ7GiKIpbN1LVjSMloWHWREVd95GOXyUtJ
Ux6RaLPGcaqnDjYgsaODOkjAZLPUcINxMKMfYSXip2WdPUgyOKolAEFn6A20qnSg6QyFGSc6Cvjf
ZkShPBThUMehk1bIYTuTRuuz+pc4VXwHXbthdfGvN6XoINZh0RXHaF1eYH9csJwvX1zXg2vj3i8l
bdV9aG0lZIYvMGZttpU+m9ejs6kpz6QxjWeQXoqmafY5nl242zEGWgyqa87cS7uIDTkdqJ70ycD/
WYURYPsGobbwSYoJALXibFzKnjDFOu4wy+3+1k5NVhRJd6zUbeB8M+pt9Uj3d9+KhcJKv6YzT00i
UCIMaIUT6iYtN9OVpJlyC3IeZuh/PsdFE1YQsM0tJfpcQiLFvjHsZmu93o1kngZDGlNkm8ygbXRl
unK7/vrPqotglrwEeFmAOc7+H6j7AC/4qQ2zx1eLHvLByQ25QEKnCjy5JRkq1u2cdTPRf2LlXkQU
mbcu7wX0vuXdqTJ0+z13e8L2vpIIjB2UbfkHYCgf//iT/S0nWrQq7edupS8gSITX3U3SItPdlJ2/
pOjBpPGhngsVxZRg8QPqtUo3QjggNTGnXxDMuYIDsF7Uw4MMpoyYKStXBnO5pxOz5jyOJJxXre90
bWf7OLKxuw0wKlKp+L+bP9eDzVQII0/J3rOn2zubzUv8HGpnflHMZZfT6k9hwXoECWT4AMupREwa
xdhuf6QGh1M+8CLzZoPr19eO+No8bKRNtpS5BW1FuU99WP9CEY9HEY6a07xCurDBqCZUJf9eluTG
9RHxewQMSVAQp8RSdBpJ+3qPTvYAkn/980hcmBV+Dv25zIvNKdpnaz9ndNyAg47U3oDNmiXhDrxz
zYM4gsHL5SoOiwe6/QLmw4hLMeJj09VJFzOtqzdkecE7OuFLF8DQovxeZX4d3+kpICat2mAb3/tb
uxOUqsfIlSUaWN/BGgL1f6oO0acnwVtnUr9OromWDhLmZlxs+fA/Ocp8P+MGsdcdzJ9lnKRY1eSb
GAlYmzGouuIdBs3odvZH6No1rr9R9vZ8WuXGCzNGEeMaD0KUPwLnv7PZwpNeUrKCDhO0C72PVk+W
lXulsuzUEKxIq0UYrjytX4yEKvYGRzXvsceVTBxc2cb5Tn2+fNSfXqwEI+jB6YSkh0SHfNYvgrU7
F5JaGiUwm4RKaYfYH8f45f5BH24PvodhUAqNyX75VJqBmP5Z+ER+zL/LR5d5LWC773wCiYfNZIi8
Ub0i4Wmu3RlvPNYyaqeCgc3AThO5NHtxmjXw+P5ljuFGr7SkfxVzCY5yB0jJZpkJNDfc0eQCX6SP
disCRnM1K+GkG1n0rQkctVfzF+tu8/uIhw7I352FfTJlWwXFFv2CIvCJani6axKtOXdpPImJ1N/6
r3jdf3vNj7DSqiC9x4SDW9D6YUvHmbptwE+q10e13tFDRo4125n9sYYTfIoZKvnBgTJ9IMCLKc8a
EQ91gbgEHVbxFGWL7Kx5YOiLEILteBy3hA0vVekoZHoL23JC03Gk/j48+AidDBH6tBHCAwG+bBOT
N7ueH0l9bhu/+ANYC9q7Lw9aaMEDMGhhDdWItIaSLVetXhYrsTaYfQTsnWUisUopV3jk5cWhiQwa
OPQVuaD35/fon1EWwHgnvHgQbVooaspHv7PObh87NVTxW2Xgg3tyrUEDlNP3vWK12QOC0ipGOcEo
MqAcR9wXkCfdT17wMmqpnmFt0/RHgfqW513RTnCcZMQp0Fd3bz9fPGt1e6lG/lOSE2nptH+JTCSg
gUyEzjrTo8xibmqqyc7vs5DHCNeCJ6RisT6SU+mmDAf1pA4nCPz8qpD50bgKxy4q4hBHgKNxNfd0
2i1J1wGCKj5/2+jVlWnt28PW7B1LoDa+KRycmhzvLVrBqX3/xOiBF6Mwd15fyoqLEPEFExtnmTAb
fma85LiqEOC8KocuPTysxYuTYuFomDTqXDei/kkx3hlLqId/v3v0GktGti/1zEdrlvSMpRbeGnHS
t6yRh90GePwxcxPZTlbMs/aWR/3hPIoq346wf7uByh2FttoWPN8ajVI+i+vLrcIU7xiJb1BJPfyl
7sNVmCXRuYjgp82uwL6qjbtuyTMNy3gP+gDbMgQ932iSHmHT8X8oNlANWCzbsQghf7RbuAxtdSI5
tCzHntl8GZ5B1Zmzfom/9N2odK5TUK6X3e3mwLsG5aayIb0aQRH8daUygNRC3Slx/isv45gdzphE
Dij3tJbp9KLn/XYg5Vn+Y3iP/aNP+VozG2rBF8qDXVRamoJtm1DiZhsL/fWFEWAQQrl7Zd2RNyN8
Ps86yJSJPh+EifhEHwQidd/VEQ/lR/zRoFTtoQF7261RAhKkPytNJneqgS9HxBVPHNYjMGseJYi4
SCDPoRMWHHHqIdowfx42B6cWHPBqqRZUQmJwJStg+tic1VoYZjMlL281nBMvXjBArL8eHWQYygpj
b1kBPK0/pNNNqGKrc3OJJNWnhgCAW9D1i2Bxq3In2szE3ZJ8Uu4ijzab64PwSgzYisWsdZuaLVIW
ceEYgZ3z93aUqfY0J0e/xWa8GoRJ58YMuXCqq4EjMdiNtTXucMV4dInmyvCVsEZY303+9JmuNrbs
/hfls9ByYk729k3cHHNgrMiMg1y9q+FlTXdLHKMosv0wrN/ptLhm+YLYQPNJvme6N8NM67n02i53
NU7MuokpfTxWiGcLzTZAsY9Rs/bU7um2MRMDL8fs5pUM35qOlUljDPUQnNo3v/+RE7uWLRJpu/cC
zsMtwmvzxM01rbtHWOoCvoh0mn+tDFB7/Pbq8coHn9pNFPOTV/gMyGL4+OY5SxD0y/6Golafn+Yf
2yr1D4UUNm2w1gJYLqZveVIef0iDOlh2yZz0a6SPiK53QYsElZcQ54nxIDwOkuQTsEBIkZhKZn0V
IfxUykKOY6KSzJiB5H+U8flmTAZR/TjmzKx10h15f0JevxrUoiqHnIDqiVgo4gye6FGbq8nmXaKN
FgrYik5713R6bw5srihaSFByC1MF/YNMsTUmdsoiXJ4qaQKsaN5/q265FfEUgOHHg0nNhDwWKfrP
epAv3/6MuVNyusK7f5+XHAfnDJpBqwfmaV8dY35nzL6fyxGONTfpfuAyLHbQH6ayIgdYLTqC22rs
yYEQEH83IorfXaYiYjn5B+bUcp38e1GZFe6FgGWHh1W1ouP86P/BqYy54cBZBSe1MwmpFy/lQ04C
KatVDXu9u4Por8J6VvPiFZbYXeJKEKrr/RhbE1N5Q9PvhnxYmYblfqcA9DRZk8+LFdNkUR+4PQfm
2UrmplVnzlN/YJnPpswJnfC6pQpkBWvSFBxCPgxC6YKezwXzF6cViQ85Ck6wTzNGuRwZJpa2zhB5
kEY2P2U1grAzxlRYxqI17yWcQzwNcLthxjc8xn+YU217UbbPkQRFmhOFxhhE03TEcFeMfZ91yNKg
Kpria/nL3bKoPf9eBXBtZQI4mkuH3Z6Wzsr+YDLtTdlHzhvA6OR151KJ9XSHpbv5OWphBx7V0aJ/
WqmQ9cpJQct2L5ZvkIvJoaxzoKCH9cUSiPZmU70T5Bu3Kuu3xCxgEjaiYjIB39vx63UzDxe6gYuz
z4mO8D2alPpjhsOAsmFxH4LKHYpQp1sLwsxs9WMaC2khbbiIWZRTOQ1Pu4fzBlsVsG3zXhohlWMc
K05dd6vF1fplXGD1qgGOv9gA1znZYUtiDmr54dKVMr29BUYTu9EqVJhOBujaR/LZNyVVlDFP71rf
eTkTuU2uozTWyQBRdrOPdT5S29HkUObWJ6d6VO3+sI4lNOR1qUmtwz0JK0rVf0uTaTteMSmVADKI
INl7FlPDF+7JqfLIiDGaBj5H7LXTTvPxICLZUOjqC1jmeaTvUaK6QpD0BUj0zXQFLCSVr+dBd6jj
rbS9zIzl7UovHd7SvAxIme4ADOFL+7Azq0jacAcE3Hs00r/E+BqsubgFLd3hzxQe5GCsHjKKWVJ1
VvxK4ext9SIoDXgsgy3FgVMzbCPvd1aCC9H/2DpTjmzimVChzTHtvyZ1CEqj/KgP3tgXGZXhwFVr
rA4WS0xqr/hZuh7xKPiK2lFYw28GlmbmOd+9WvZnT5N7CiG2STOMdDTxCZOV4s7pcVF/XfeU196s
8zyJ7DtNxLuqhhpbCYEwUkQfyfBjTpHNripY0I9zNlUTXCXdJtvpeQ8jnnpoSD6Jl4voC0ysxqik
Otyj3nbxQSBcFvKH9ATu0n9DCqx/zGzgoOTsyXOjchwIbLeFJlafh+FoeqtJP5xqV4rWSJ7V9Ma4
2v0PCqYeLiKXX1pkWNVue6MRjMDolQmM0Q/Ac9kGilDnAIYNfYNKWRrMGHjIc5/UC+W7v1/Vg3Pw
jbDdh9cvDoAx/C3RzfBsdam0q7UiKi+hs0Jz+NpNe1t86iReeMdOLYhobiwwAiyD8PoHdN67d1dL
XG+HFxZxSC2uAd39RHoCuSN3CtlnOze2SmuSmajB1BZ8lbyt1p5gKDcghSMCTdCvArUVsvUQJCxX
5fk9DKvH5YbARxOoRZ6w/Xu39tuUlCrxNz2n/kijiBZDU512eyQeOnFAfBTuNraqYbUWw+HkqdYS
w7BaY/Ns1/nrBubYSFZ7+sMlbn4UHuu4wYs70QJiCPKVMRkjS57YlT1CPp4jS3jcWqptBtxGBZEA
Pa7h56xVHh4mapCTVnB/KtanbN1QjQz9YgP0T2sXLJhMeV+Pdgg21sEew6Q+KOs3f+KhILiZQLQN
prcThPitU0aSuI/NU9vogkDwUy6MxvlHOg6zG093FfDrSdcxqfgurT4XooYtYVfKrfia8ATvDQ0z
24fkqLmnlkRRLI99YEqyzI42iwnlRGf35lCdPCoR49LO35KzqUCgVm+kc2nV6Ji/GxbYTSTnXe26
eHnjPZ+dmU9B3VZWA6FbDoy2fAZ26BrOdKOmXgcChE50LauoCiLFMZqw6LqmJ8jMtjV4xvWEgozW
0nIBT0ZDnI7meUtAic5SC3fZg/jG+LeogOVV8SiP39aIDIurRzIKRzNXOoBRvounclXpJHYPONKt
62JmPbycPcvFzZ7jZxXWF9DghWrkuINRgVUcCbPgXo5v0hWXSg1et9unXvKqoVoVCxKgDtljWugM
GZMj2gGEZaEbSYp+WB8teHxVN5kTO3uG2VUApNB6WOoOKwSoMzAUKq7ctB7laptMi7hvoaHd1m2T
Bkpx6L6fiUwSlwALSoRQq9XR8QynPIysLVxUvZJ+Xme+/m8l4BI50szVIamv7dZJpef1JUfRRGgl
vjtr8DkFB86D34+87q6SY2HE8HIHD7+vu4JsZIqiJvHZLyCWtYQRksrsIJ7xBBrvLd8UVHp1wZlp
gdIRUL5sybeGyI3q9DpkyvBDo0ha6NV9GUhy8T/v1MgTaP04koWZ295rvKepF5poSesxkGoubz2m
zyyxz02ciTZ4X+aSQqk8pTVZwWyC7D5bFrmK7lgktvjxy255Ua8SsZ1ihIUXQjnQhql8KH8f04i7
NeezV135/m4m67AhvErI7/K3099u3Wz/s6qdffJ2oV+2TSFAfh4/1iQaJqxeZWtT8lJF1gDMGCeJ
ire6iu3tYkEG3CRxieMddkMpSSHLMLRWYr6wCJTlATuBaa5Y7gGkZejPJ0jER3bsK9U6C/ROIqhI
didS5+qif1iNWh2hD91H09mzGTboPTXBlajss6hq9lUaUBZaw/I4icHsec/KDQYWsdokiPb3SvKH
QTQ88v6Xcb0eUbpN2TOJMCL+cWFtJDbaoCoMpG+NLKsFaWxnrcpqv1Ecm2nS5kb5fnUdPszC8Po3
J3yO98fnm4j1sPQHPfEycptqS6LYD4Vk4a1cGlAx4FxSogdcMBUf6cF0L2CXyRLz/bvUatTg/pPw
ctoMfKSz+bxYEHpgKxV63/U3WU9ozrZjT4b6bajJ6ru6wZuWGOj4vjEGxmp52yxHNbqFlVecJSvJ
nXhYjYr4h6S667fJqzAS4k2pxwOp14OH/ySr5XuxRly9zt21Szi9eD4eWWSigac6O2yV+VvYVkx+
KIOORQK7iiPsPwNOaIgxw0ykvaXNMJmFVm7cCPZ9t5N0P7MTj+euo9h/Slpvk3oh4dlWp3b4oaCn
vWqYq79eUCxTGfcj0Yc6YL1eqPvYF5BD8nAdHvUzpAZUXhNSPY3S4RBjjyq8+yBiCE1FS1gx3FPA
1xjE1/T+fgCFkly0MwDZeYL40Hq9bASWTEGSaPQ1JSv0ektd1bfMus2E5nl0FG84B/oGfOZ+4+r5
QjjkIB18rNazcsNyR7cYDNwDNivZgjDF/tZkNFjHywm3ndOfxSSoNyJjeNIxULpjXJPzVzQuXrWe
gQmfEpn+lYp68AVT+04jTVZRkdD8Y+dXNjKpQ3KPRapvS9lAtdQDFbVO9B6vPBoEadZSO7srgnD7
on/fRQgb6UWic/bx3wwxsCXCssxZuX5Wb+pvcRfc4sL2CkvRiZyS54qyn2oGFTPKplxY3J8LQB4y
dXDjjwXiAVuIc/MMzdYkCpdloc+6BbWSrSdDQgq2TfA3W8ZpTMFiJTaMswvLpxPROgDoDLGVeFeD
ykLdPZnPEwy1R0qhQnFcbMsLXSoJK6C0LNzKe73G7rDcQzkrosx85bg9nwwijQ/pYFYn6fYUrvsX
7E4eTn2UtZTeKaGXcaIQAXHQHiY/eC3pfKibphzrYE3rv5z7czUEIuZdHFLcvTlLRpl7X6VXC3Fi
DBSAZkjJb08WRAVhzYtrqf/3XR3ESJteWMg++wG+WCxQzxcneSIdsIPxlmOuzd291w6rhZKXhvOA
hipXBeopj5i+ybSwLkd4dF/c0itBPjmhSC0yxsHvmycsokc3eFfGyT8w2w08aqlf/hh42q8UZpEq
J6j7Lh4dtniNSQ4UanbrEEnw9+ZmbJlE9iI8pdbUhYpyltjDKZjuIbNk3nAvscc79zvWbzXFx2js
YVMCGRl5KrlHtEaJ7Fg96h71Z4M835dbUqoZv2bA6gD38wyd6xbLdFL951CrksN3nDmCVUDY6oAv
p1BfbPl3BJwfcdUQuZAIlj1jAEgaU1RdweMJRQpZT+uLjcPqWr3/IrBE4AMk0ND4O8FmqwuPecSP
anCobQw6oxP4oQQ5t4UY5o/LPe8qHqn77oSezaINy5nBFh/R4caZv6KT/9TR0+uErw/ku/GOd8wV
ttveHC/rHu2Z2WYgIR42239w2h6lULhsWO3L3SkSb9mJ75B08UWtWTBuFDTjSjBXECCBm4BZHCMN
Lp3ms3O5or+UpPbeCMIa66ypGqHKIIV92r3ReZXhxdYCZGVK1Ykzz7l736RUo5yF4ywe7k6rWwTO
7pxsE13QQZSNXjIe5OTvm7K0MjzSbJ7QhfiFb+9r3ysb4NbIxeU8N6bo7CQHZMGcOzJy2ubr5mbM
1yFCEJMgfxR3256MIAzzj3MjXs4w3M9Omg+PkaL56IlrpgX0XyXKRQMvR56hq85Bb/soMhTvluUb
fxDTdYCjx56p3AbfLp5XJumFGXQywWnubls5GXxSBZbLzmFlvpN7O3C/I+dTw0QiQC99UQEV+VXW
Dy8MTEe2crcG1DkUHOhilMD5Cs73H/2lslyIDr8E9PExo7qKahEVhNSzNp87Si3MalqmmEfYCsfV
lm4tT9IDggxoUo1sUXhI5ozNe7bpHtkmGU8bO4ccaaAi12IYEGNhOhe/1cphdd+dx14DMwPVjGcu
44iTvyw1/J5gnSAPBop+LJJi/RRn1CfPYae5n6w7LobGHHrqgxQK17bV2VdeKMmyIzy7jMQG9ZUe
RN3+y40n7z7bUvvKiEDgJRgliO+mWYbMSXt1APaSXSkdN6/0xgp96mH3J0Tz+a3qHaG5ZmThI6j2
QRiy5DW0ziaQk9h6E/43oURlS3ieduG/oeYDHZr4DTX2fM4TjrbWWwneDNSOuR7PBQxHCAyaCxTq
KTqFv3+AsEU9fYeT/CpkzdaU5oZpXdelDzbZM/t6pWwgURyFsTI9cqE06wuwAYBzq1Rr68gJGTX/
eDHN4G4m8ZIfygkF0ui3TJ2NmKQcil6OS4FGLv0jJZgiUE68kA5+1ZJPJBQWRINNd8i+AG4sWGPi
fsMtJascZa32urwMofNzY6P5UEKMWPFppm17w7C+zW1iqZTi1bYWOuDsXvBlpuWYAYEa3Z9qfpaV
MfIBfnxNJgmV3IlOEsEXg23LD40odCYQRCLPmbA2UWialIIQ/ybA/B7ZBjmsl91O0X4FG3jGVJJp
u6KOlSGTYItR8Q0pY4n6V2y715DUdf2iEk1lHgu7ShroJeN8MZlXPkI12qHfdIz22salceYl/qYQ
2nbz8uJCUWViwsMY3h/VjN+HhYSkuuAPzaPTUMLoBMqqqgvdinkeH25XyrJAj4cKFfCIKexktrsL
mM9f+RqRKE34CdNhznBMOfcNFfIpTSCAoklHOB5XP5SvR+4y/thiCsmkopKGiiSEo9xD6gvSYHZZ
uPDBPV+JdQIQt+QX8nYXLE1G1ELyVInSXfLrg67fS1kzUxP8WAop6KGK2JNwnacPZEQN7hNvs489
UZTWuKKnJLr90K8HbMyiRcAWIq0GekqgFE+QXEiIfq+afzR7le1Cr6DsXVKgo1GIJgNEp4xeUGlS
b6XV+UMJA1/014PJCGoRnmoPqpUiR+bIaFvjqQW4AKOHHqsYif32K2iMuD3w4f3NfQ2BLqNquRJi
xzNakPTeydbP+TqRu28++bUdOLnaabQjMUXRP/aQ6lDP5y0fdfB/7pSdpSXxT14t+Q4GdHQymL8l
Bg8F5TMYikJfVBAypnezAEFLNC3y/DU8tvx6kZse/Bcwtm+G/RoqDdLxGfpd2TvuwHb1vJkblsAx
sGeEr7JthSBXuyoPk5MkaIh5h8yljb/Y6ptuTE1IP2wq40UZpk2Gy9wn5UqcMDVcW9SiE2UDs4ye
4VWE90i4JlKCB+yJibF898NAYH6DHV5idDBr7unFoRHyGcy/Fmed/U7MqBTZGanKgzqbsdA+KwSw
PIEhhDmzusSU+iiiyM8GrRXAFW7n7I3o7p/QUG+tuCP2SRwH2MtGPe7asRbdyICOdx7IDSCJHGv+
TCPEt+Yy4vkeMs6I2kZ+8gzap9lI7rjkK3UZ67alTwNMu6KA8bq6L17TpCHzQw5i8/n9NZGvIcpp
JTH0fBfCiCPjDvt54JCQhu9wkjFTmcSM9c8ysjJWCjmgbvJ8jh1A0ri8SRj+7l4BQSjn2Vlu1lPO
axnRHyaFDrFFNvQximdzd+J796xHEZndw/lSc918Ov8niXuaKBaa+lAnT/n0IgDUauVOjfBVUDYt
gjDbLAFdYggXqnOENfFQShG7TDRn/Po4PkMYZR41FqIHsQoGr0VbCy5rIqODAjfdrBQeeCLJOMcC
DbRqRwyvBM5eOBmdZSH/i9V6De7qV3QORWSADDOQj9grfv7wXCgL4H8++f/0ZFY07nt8PPkKam57
E6Vaqcq76YLLSZqxkXjVDKs2CdlZPQ/D5oyZF6J29V9antgFlcoEbaZXJqXDGnf7J62UWjyJMFTh
VzBCW7KNt0Pih70swOSPziTDr3SuQlgJ7OUtkJdUkMHnUDox/Rw6v6IzXfGAaq4EqLXBA8DYJYcz
L6w6CHzlKtui69wplravj/m3YctkmgXTZ1pDRsFrHMfOa3QJyuPDIEs5Rl7KHTcw48jo54x4ZaaP
1T5K0+T4tPrVnOdOEhZhc8qLDwX2Q45aj5ULazuPEtbj/2naKEBcpnz/EDaXt+5hbYHdfnGPZPXC
o29CrZVGDcv1Km9lFE1qpccFsyQmwUSkHAjgdQeazQH25hxqQjOoftGPTvsKQgxUjN3DM1JNdZeq
rK0uuannizjGSZD2EEZ7nHVHbGMVR1390nm9A7LY8NNKef5n/KsjBF9bgwRe9zuHWrh7uQLTu1XA
KMl8q3h2ECuE3LCyXhz9zkfwb8357ayUNNxDl86fZJrXFvowm9o6oqqkV2rzI/UwG4SW6UIBL/Kq
nXk1VjN9Ffn1qJCJZhv2cOwo5m9VXzE23gKpB6ofP7VXMoDAqJj1Q9eey/ydtak656WcCN7WIlJ+
Qf4LdbgijdTNg/9stG4qy3kNkgsbWqPaDhzFFeD9aKsEhSLDkmeGMc6GtT604xfFV020P9GJ/nrV
/Ryph13KF8TTzlOny8OMNVr4nP21AxQh0wBgp3uPUxjN5cKjIcGJ78IrDk1E+A/VbGwwEcCVZ1bh
tS7DVk9NZ9HfoZhwRNVWOyDXtgO3GjOw4YpwOWCvk7iahJ/1gDnbUnKerHTGFxF9TmXqYaLD/lIQ
y1sYDOHHLk9LYOu8jgEbyU+2zhKm+Lf3RvC2kgwyJPbCnQ4cy83mzpHaSuUjEvNCMRz/FH72sHdQ
ivQLw2HwcUUPnqO+mf0nBDupXnKiRxqTonl3g7zJlqzjnnXAQ4mfl56jxOvBMkXVaUNccaB2MH/x
lLrlrCzyyZHrhZJ9Sn4QoM249Xzz+lZISIpxCiQ4BEpiDPEf+aafuOLSqhgTZch9jaXStV1EiWPr
qS4Aw1PuxysvPVBxO8rq559bBtb+2oY0J7qxaw+LgLK4FhdEJZZKMWYqLQwcx02bk2QMEyImTjaA
NO2uHuqNdZ2p2nSTC0N02ytUnPEK9b+9iZCQ+Zy2eyTvE4YJCEXzVqx2Z3XZX7153HF7W31nKumd
NeHSw+Gjk4hgiINxKnZ02bx7YLBhNF9TVluyv4plq1+yE0O15wulQnEQmOin1BC5j5+wKE3UeEwF
e8wMx9n4iboRNzOqaL/bqQyoq5gqlt2U8v/KBvOMQ0Vsuu7mmctMvbXghlyk6LQ6hfGnhsFnWYn1
vIbaRXpeGddst4n/gCrs+O21eII/LKrFvnVSyZ4xPOTBahLtHo8E1cwuTrJMI8leNjD6mT2BHrLB
E1zQCLSijeka2z99jKeTIyl69E1T/b6TfeH7ow0K/IMvyaejevcN5sa/CK0dXtduLGAHQb+aWtFi
uI71J73rKN/jOHFTYwVgy738ifzbHWdoimzkRYVwnxG4DcuV1EO6jcmviisGuU3mHSShvh6Jq5bb
HBJakA/Re3qlnLnnVlRRY2/i7zG7tXO0PJJP/7MHTNsxmTvvS0YUPXfP1wzsRvGflskvTCgKEFSa
kxjFGCFzpTuMpyOXiv3oh3/ZDGqoS2W+du0rYtBeooNYk7eAzlluXaZiqZV5Mgks3jfUXxnYWKiK
2klYWGJ8NAlXmygmOEh3lDHMyUcRBpQRR5+lyroI95VHocMAozXfTYn0Ef1ZHrvKlob7YlF5kvIi
opC6dMQ2swIbH2GNYeikY92v0fcre1UG5QQDIg5le8h3GSm9Ujy3NtyQnmoWcAuTScNi3dgNKA+l
Bq3tPOF4uZKwr3xQvNS3+IDaHCG41zna6Es9Q1jma23eTqRBEK61ZHXKQZ8++Fm1neIXdHN0gvln
Yv5cvPPPS95blYkMuD8JjhPZi9YQ+/1Mm+2o1UJPVuqhD0Owx/jW2MZTafodDYA9mdrkElSQyrMQ
Kr/KS6SAPTcrYZBL8cK+r0ZuTpxt33jaeQvqfNASpE4zmdAR+PJ69p6MvAUCCr5V1bLRZhjWAQ14
JPcJw//PzmxOLF8cYgYw8pIa0yM2OY+DM3LVkvhN5FW7E9QqJVqFvRWgIYSjxfhVxWwWK4xAmQVJ
803IuX8zVrudwQuhjapyeGiCqzXiWbPyaSVd54xWm+vtSLn11MW8Doo5fokKFLuiRT9JyP/8OEbK
uyTYjCKxWWwok/8lRm2DDywoQ215P1aqZD3aSYTzIvXj+5Os1vSjbxI0dOQw+QHfpnXfhkQnc1jE
k1WZsgSeZpqiQZCITzuQ42JKEhhUgKYd5kc2kaKCJIN2Nt+b4mQ8ToJLfZkSjbVRtc1S18BvWP8S
U7E10ulmd0ixN0rLhIv7UHC65VWIOKvpLXs+mUYTiMSnV+6IUNr2fKC0uKXPtyfISup/ohI7TpU1
qa7kMynCmFgJNTFYxDvffIYzuy2wEt0cv23tFCoMCGDFzNsptkS+ImbE6B0DYmA0y314a470YJQJ
OcvBl2tMK+Yubrc53FZs7ls2jamk3GOWQVCE2ZyOb/UGGe03W3eGxCoSlqmAlPNscBkGGaiAITOg
4i/nmZ1jHiKb82xmtBmSh4hw4cZet/uqI8zeoCm306/4P2eHd7o6EP3JUgH21SwuOPhvmY7tUl5d
DMv1zAInydrZfhVNg9CZ0SNW19oYZN/T8Z0HKuPPmJevXExckVLwCb+H5XBgzTlq7QS1Q4qZ2p7K
tQYJf9NLyu9VIBt4oAqgpBvOq3WSqztT9zNqFhrUSztz7jSYVoMSNTwxLXtmWTuTXaQMYR5zmNd3
Crca46fbbqL5TjbQY7IdmE9m/A4yNRzsgJn/9wx/WcCIZL8qsVmVZMhyeuaK9OBwk4v1cTNHPAIm
uSHSD2pz6izxqHWrRchdsUis7cjE1ybSLOYuduHCdLgleri7Vy9DZg/K2vpZJnKaKg0PpqeC2YO/
PTDxcUBPNAuIsDCQN7T/bO29Np64a1sbWatbnR5pn698tPylT0FvR1DOEMHdAqArBQkeZ4Lox7nf
qLMokmaNa3qPDKTHTQDBpJUQsWnwXGZnmILrF4enLN1ioFuozdN39a307/qKI5gFSCvwP9FB2L1b
awL1Soa2wNQ7wY6dOTZvXAStfa2nmMtMi4N3/W8nymh4xreZEAmh9Nh9gSy3jlWd3PAVTGqpN8Sw
ZexE7vBdutcpslwoYVVc7Cd5YbH0d815s+Q87zvO1UDLZPLpXEUo6F3MaQNsHIO1xcv0esSU6RX3
LFlef/B9ccgLMEUpjC5SkpeERrOLNJ13c5bJ5zS0UY3mL33TSyKQlqPSmfZ8iQ77rih8GKKWyd5K
atsaIURXlOFq72jRTCyQBe/Yx6KJJ2p2onxHSmZtapNculWeU657hdOGCu4P/4f4mv4pyOaUSQys
E1riqziI+u31CrniMw5dSmOj3cZ+dZGanG5KPqxzoi+wCz1iNepOPMOfd8R19C2whQi9h0SAmZFX
NBf1ciwJeeZWEBxsK8AV+1dJzcEjBbXOmIShbBC4BU1JYmHuFPT91AxUlZG0XeDqacl/lIA4rO4d
lyXGVRR5dzKQy4SfsGivT34hjyEwyA+Qj8WFiTtVn9RejGnHCbHPzAaC1vehQ804fVHFBy0bRea/
mWuoONtEUsfVVXf+sDplGacB26qrAqmHCFsO4XCD5Vfskl1IqkvpenHzTiEnTKWhlx78AyBlw8LT
hLLeJVJ9r4Qj2XGdJ4PZ+s10uKI1BNPT0ZLRiceg+grHeWzSKdVZBgD+S9ZE6nYSri7g/abUIgKd
eW4uAAQRkzUJs8OJ8WQDk6mS+zZgKDFk8TH1Em21dXTHn3v84Rqhrm3KI88orceyRAXGTEhkVfki
a7kfH3gLws7kYR+lFVdtQ30O11Zh7VVpTdcOe7C5Dx5bcC9TDKmH8isNWi9nOdD1vEmp2LEiwQhb
Fhf+8aFAEx3n6+ioRKle7wm3S2i4N9qBoTMxvDNu+ncPhq/9LiXYBqYvM70Gsq5Gp1GEQpRajfxi
31LBZJAiYspQrWK3CLqgxKVLJKZ2G6cbrDTEsJL2mAlSX6gaLd4HVToQPATtI3han20Iwii31/J3
8oGCUwwrBsTvMYlpl/xKe8JG9Pucr4OvDKxHXnrOPun6wLNpO0PIIbd/6+RpfiH50717lj4rtRiE
3Hfu4fASpeExIGWyhBWkQMBlkiwokVeFXbVMwIMkMfpDfFp2gkTF6rXvD1/rKfiuJo8yaOJOBm/6
II8fuP7Qh+yY/FssHqaCt0kszGfYUNxPTDnJgPrFItK+Lp118qM6WZQRWuMbIX0pNhTE75p4d8a9
6be0c9/Bjxhu7ppL+TmzFZFiOv6wHVeJYpHaSpiGigElwvtb2cUR59enyOTqtpqXzDKOotBID73f
gDM8G1JjRPLRaZynZLnae6yxTl74UW4o4iaTQBB7c7CWjjAFSt2pF15Ertg5YMzPe+MdePPbuiYg
mtMKcljjEerPCEhQemwU/M33jL3SR4wg4rNbPbSBi8EhvK3mVR0GZfZDOZVgM+ich2t3mQEJqu3X
eb3hieIbxEsCBUy0ir5u3i9EpKMZroW+V4yS5i76bhd2uGuhPJnGskAANDNwvPIBfZ+NOLDfvqVQ
cZn7tH3bz54hNnLXC9q8Dh5jK7Utdu+jtNg268+gRmcG9JV/OZbVIfO6oR+T6AfJl+3/dVc2iCV5
d34y8Qm8+jpKoErr2CGESHPpp30op/URrLCHSVhK8J317Yec2ruumml/RuytCAxvCnPYpKO2pvDx
v/v+mnwawtSt4ckXFOCulYHkEQ0UNAGG9jEhYoUAjKmFThp6A6zHNhsqzn0eISIyWAXObfk3s0Z8
Pt+ata6HMKqDZ4vfmGe1m0d6YTcBQv31oyEZjaaPitAB/yIOC/4Ptzm7315vyW0Ls8lR0ohvnmEb
Nil2aeuAxdaDK952WQtFGYlMv3drLtzeGIOX5P9FSC17o1qz59VchRj054QE49WRATYss9nA0dpm
kJfUK1PurHw4z0rHp+5doj5iSTTv2aGCmhid7nd+raVFoK96KGtwUDgHfIx6OWLGYn0iO7Pdi4Ve
5aLoImbUvy8r6JDr18BH3HsriiL+AnkatV8je2rBXbh9GiPIGfrVvz5qWhvo2RgGukZLiQJabdji
L4Entz2j+QhDPWe4QyhmC8Ci8nxZhSIUWMbOhpWXwIdySjwsv5xiKP6X6VP+OMj9O6IQnjztWATJ
PJofkvo1IwFTLuy9OVTKAxRPrkdWzLac0VlQEn5MVimzSQAtNsTu8Sl5l6jnCESfuQ4gzCqygwT3
a8g7lh/TreVOoK9R3WRD+1UCYODT0naf5/07PRmNd24ZKbdJmX39YuLF/Dna4NhBcq5woECJFi9/
igmyxR0o2fl0oI0P5dJTtuOtbtcfqFG5gwkl9d31m7gyODNymjLmg7sCBA9ECCcgBAVyJ6x7D7XV
7e/Ov9I4OYs4zD5L7t8pDSS6Zt14pJqsjJDdznE8Ek15/HTwSdvGkxeZkZnD/ikgtlH51gnPWwhg
PuNIvqvNX9wcbGHxQCqLaUubfkkuJ8pRsxB6hsDH+lJgM3ouHStHlmh1w619yAyGyZJelUymQmrR
7E5qpV0b9cC3ozZTO4NlUJBuiXi9Lqd4CPYDoL5wqQ5VeWAs6CoCUmyLrgAGZBaYLzLXZCF4DRUi
HypdiqeIj/YxyATEltkk0KLAFVqM3G1KGCST5t74rfMoFKzkaUpcpvJhHmRwXtiDNCFOsfaYG2au
/RVrIOl6Fd+M30anUwBV4XBDFkwpYSFFv4ZKKq2Kdg6bOus4EVN8dEKC5W9bokmceWBok8hf+mel
H6lsTmNwVp411YH7A8uS0TnbQiKlaHRxOlLYjHao7cUjcNGjeIl/3WxFBXaZREo95xdQlnv2GIZj
TashDW6bwbsFwUi2yGcEK90q3uecoOTH7G60Olr+i+AySaf2X5243+HHd2P93h15e+ZeAn7dSOhO
rr31QKGd145qU2uug/PWpUVzz0Fa5CCWMPJNNoQKNXbnw5xbZmlBAjOwexNnoKzO1Sg3d/PKFID+
aprAoY/QFR2cWHKA8u+VjC29ZJfZCuQZrVBHBjedAoJgW0XEKEa97MJpDxXw+SyksHUuwAsU1FY5
yTHEmW1WxCn/tqU0IQcKuBnmD4sFsJpsP6LRjSc2buyJKK7gNgKRH8em+t6zB03szNeRhH0r4P2l
c28lwFrkWKZR54OWCl+nPjR5bZRS42YhcZrImAXrDcCg47BSj2uMQPvr+X95yla7EdhCplZJrdAp
+BguWnYzyfv5WQmHoxp8G8XdwP9GZXPQjuhxTd2DrHIDmfVm+pStGa7sv3JGqhCVJkOJocpEO3B4
6TuZUbQ0h5sIyZdMdusXfPsiCa57bqqEqYG3E4N86WYB6anIHZyIQV/R14+gQx7XTY2O+z7exJq4
nX9t/6y5/VomxHsSYdl9y3fQ8LvT19UmjiF9LMPlY6csYmfByNilEgV/dr7CEukpMYdgXcu/53Z3
0a0ahfXlW0MTiFCWfLag5ATzFCZNVlHeFSSBt22GgGkizvYXD8KGYYkSKV1NuDkxtAnv90sZIcxH
OtpUqiWeRCz42ugDjSQbgS2/egC6BLFx+/XUIAKeNP02aIPGX8qVcoBS6zE3iCHApnyE2p337f08
xP1hkBMz0dohW54Kr3HO+FOioz9lgX24XmySmpXc37P+HbnZs0NE7uCEexU3oShXyE/nLMWb3aw+
z4vC5BIL4b2XVJLv5/TaqdHbH0/d9SbSlLr8s3P58Q5Ra3R/KLrNaujDYZ0gv4+1WC840vZiZzjd
2NEI65lHyXEuS+ZmLXCYwwIciGZIyssZIVim/CVXU2jmmH/QDOQ8UpwWoNgGbLsWMl2NnoOCjWn7
cf+adLJozIkl9q7PyecuVWlZUX46dLbDjarDLbEbEUCMObL1oOkX5HWopxC7xtJE0S0767EBj5Jq
4zljT2fZlPJkRZVgfX0lAHN62fH0RSi2E5RrkXiz7YjUrZ/FZXjXi2I899h+tY1jIvd4wheNB3uP
UwCj9h7enBa+2Rgv17XxgEb5a1YYz6d+9UyN72c/5Y0Nv0FyqYr2US2o91aakwisTBCTIjqcaEr0
sX71HiwF6y+As3ANgKvQZp2uTbbiZl9Rm8NOpb39gzhiZjNGM3GGsG2H330td/uX0wxSJOznr2uo
jFhXw4RhXDP5xzmpZkB551z7IDeItjq9VYEoNYPyzTF77iWxMFO5QMSC2gxZe7gmGwATfbR/VnHz
/Sn90tkRxlyk9h8H0EO7bLZ6CcIMFxlY+1QiWNDKQgzDpd+d/e3C09J64PZgqqvHk48QUOYjmK8E
Rkw6WiET7JKLWx3x9VNlG8d/cnz8nfo0BSj/OsBzeDK2WhdVZf3ZNd/3yCnuLPADosrP6tAIOp3P
2fz48NAkuXFdKkuQOHQ5fM8PI5+PWC576wuUB8qjBvbr0SJkiajq7C7c4C3Zu1FQz507jmyNC6QC
XSyPJs8tvqwO+rmGQv/RSBgqmyRGh5qFJPQnl9g5CDRATrQsznUhjSl8+Sy4c4frk8lvAe+rSOed
DrJJSNaYa3UwTnwJg8RdLgH/waLrnZeBgZKeguPUPVqNEE8PD87Istxo6rHFp/0yZfucGHKTakNR
Jb0TmLBq7zedRZmoWRxXlL6/OoJdfozgnM3nbfujmXrZ9N2vi6ppvLCht6KZeRKvKo+v6P6OcQ9c
1s1HYYPwOTqhNHjA68voFdD4CJKHBYax6mbVSlFpvmC6jIvjMxSAI4g6pqzePvks3syOVxxlZsqU
uxQ+BGj9ZutePvI41lxVjSw62tO7R+JqliuAkfhIwYBVUfJZGpqTxwAr3y2kR5IFKbF24VDTBh7h
S0uQw4QEWN8n/QBy5P458IHssZxkzM1dC600PyGHsi5sYc74KyIO3vdgh8zKNT2uXmEVkiDpNJv5
Udc8PZCbRoPALiHbByr9MokjR2a+h5RvzT8+Tu5esxPf6Mfowz56ZZ8nRvJUkhOG2+ze069Jgh3u
khoJa7Lz05Fo561ywnUSRaTVNivYYtn5FyL2yO+8NSxMRHoEGK5cyafUXkLpHTcUfD++hG//dnB9
cdSTqK4QxPtBD0JwCGC6v/azughS4mgfXNQ6XJhLkGUDklcCqwXTtv2GnzHHXfCZ3PMuRhp5oVLu
aAC87e2da3wVhpw0tRHacmrGmyWdJC4lSoeq4BwlvIyQyTbOVOt7zP5XMspFb6awSii2BR39Wwr+
V/l1sv/JVGxiBD2YzdsxUqVxwqX7HEor0KgllRHbab+MB4SFZ1coeXG10kmUv8ALHmyfFiHO/BOn
02XGbNAeL97RSM+IS/7toOc02z3i0KM69dDcfEaW3yE3Qj1wBZZfizYhNckDdYglbDCwUOV1Ll8a
3useperasxf1cwMrQ2fDoJeyMvh7XVqGGEbRZVueiG1GWydwzBQW4+fVaR4W7DPxb3HWkQfB+tkk
aj6M5qYQ6+JuCjJC6wIke3XYmJeAo8g2/ewRZuNYAvShZ8NSVdSsVtN3FkLdsQNAkhtUpidg/8hM
0D1em8b0ozvOwCqhcDv4xqsooj50HL2BD234MADrr5Yw3MbTlFBjV7DfIVbFhvziQzUVqkDRvJS3
x4vuuuKj2J12JHapbDHTxfBJe8T08nTHZD5MYZKF9NxF8/BV0gq7pSbD7cb6nezzKPO+gTlGQ/Uc
DliVagSfH979RW0ZzJ+BCG6Kwg6usSno67E/fn5JNnUrinwzRCS0GjckdzFONPu7TvWxmXWC4rXn
5f/6RXb6Q4vJMGnRWm2wBWkxdE/cKTVIGs6FRENkkRQ7WJ19mOfD3OB4KKS+Ny54Oyp4y3x+nU09
Sfuz4pfOsz7NlfbkhZnjERNyenEit1U0KsN2UVmcUy4V3dGQwQ/fM177q9/6s469/rBT2EcdYoFU
K2DQEtspQJOq/Rkx/TkyqU7p2rgWuWljpgDB7kykaB3FsEr3O/gFAk6yLGOTBeCsdSi9Bkq6Lv9I
Dd5CF4Vr5att7WqjHnamkTX36aHy6GMU6XWd8JEyv0iz80WbUU3r5h4iFOS1wUJONjWm+cKMv7RF
rmciTOrIEACiT/90tcP2H6kkAP6Dj+t4+l9XgQscgS60fPyrtyYiMlig4BIHwhDHM+hRP8kOcrNr
5qcojephtdTlUDNgdpNzIAeezNsQGQ7H/jCcVJ8Ha6bGKe6MAmAPE5+L3V10YnsmBMNAzL3UfJm3
O+QYtfbQ7wUKAPkC6nwIElzHl6NUDqEOAYYsq5bWqnXsLnHRGQxFD+OiYoknQEgB2YlR60aQadUn
1LBX2bsGJLT0k5BaQ1tzp2Qost7jtlmtXAma4i30SM1mLwEp25OneNdbW9Kar50xEfvGhmuvzCk8
LsW7tZEFB3P3dJp4ghAOg4MELHVhyaaGur5/CPfF4dSbruThRksme8qcjfl3C7IC5q1j1tPL0ieR
d9HId39UbW9X6W6fUokfmiaFVK6UYAjG/kWvSx29dO7StnFWyhRopqar6zr0hHJpi/U/597neKsM
jXKvVCzzHRi6wPV128QGAJBvbt51ndTLuLXfHZJ80ErVkfMA0oRQDphAt741hw94lLWq6F2OIvet
FgTdbWIgEzDGQffIs/AxUiJUuJTyVl7qgHzgMA1JqL0utaJT2HCGILDKCglWMvEW72wuS1/iHm0q
Lo3z1LCFYdJ3RFJP6yq6dOvBh+vzhRUfNLxxYOWEDlZozNbNPHPFcpYiGBY41jQHxg3gI4HDZUVc
7dslCy9kIFngdLRQYriJ6JFgmEM9VbQnipPKN2QZMKJ6UrlC6UpRGrq0G4mXPpN8Hayx6a8GdPjK
4tn8XAPBv2bBqmWSKlNh2ZxaEJQ7B8geUgzrUoFYu1L0yODAhZ5xCflEE2Nfae8+2Qtm79oLGSmm
anThzo2wvyP1p/t3VtmI8mh0ZzFz04fy9yIUV39gdFeNcPBOHkxSUjk1R/vee8d1ZyuQZ6mMZuSa
2bOHnuWySnrXryquSw1TBdD7WihD8aoSyLbRAKtWJXk+od+Ia8WCcDMStCJinASM9kVkbUrb9Yba
iARrPPX34ei2b4E0eOLk7i+4wuA2W9xxfTFmJdaoAM9ChNvMFnnOtk/WoRWgMw6MReBsXujO/4fb
YjGfMCaFgt1EagtA9r4iZXswZGBFZTukH9CXUTzF4BeqSIDslJdovoqry328jpAevsuMJ2EWgI9M
T/4WbNR6/b9ind7BSUrHMPlIITQnSirNLtr4cm11r8yrbTgWM4Vz1i5D2FmuXGTVxhl+U0RKX85v
vv1iDIXTXLy0X5tJauEAytVvuQjkx9HmMAhdmHiIiQ3xh8glsdtQQ7IC8zgsUINLfWoc7ndxO01c
Zi3Vi4ylQEoW4NuSkNvTPZianXt+1sL+ntXxBE4KtfXvnd8hYbRgAAOwW0z1FBq9UrdgnIWACkBs
2bQOd8IwihZ4w+Lw1wgQwYQbt4qRE4TlKf+a/gmVYzgWG08UMXDjTyIM7qMVN4EEKmNdIYYjM+4N
vz7f1Gb8GK1MI+nNurH522TqmdWD4aTzpiQGmM8u6JMDxtOzaPtbwGv/ZlnVQMoS5Uc02KuA1s9+
iwCs/95GGOwEn1FZ6eghFrKq2s2LGmTjBhX2WwkNEFBqqml415F/L5HrnEZxuxNrNyDczeAheB0r
4Y+EG1TMvor8n+QSJWQP/d/q5fF6oj9hdccElVbDAxYDQUUHPjnvyP+AH5wYUASbCpPERWti78dD
01902aAcfZafItHHTh3CmuK2GSVG+epMLOVsRxAER6PxmEGJPYXlZHNIus/EKSG1x4BUqfVp1EsF
lgtxBqKezEaD52UtUCWV8FvVEGNCkI245d1NkJZzcf0R1jNkdny7IEmHAU3IDuHFVvqF1YRXFwQ0
Jyua9HM8lFf73EQJJoXmiYY6jqDvK+rKf/qQBMYlaNETpEnEyDFmbz0qK7O0BIyDZbQ7CAXeqpXp
mFqCU1cAYZ/egw/2ewfLnIBsa+UenO1CbSEAKth7UITRpip9xBuXwtgazP88NXBX68RbMsUQXI0u
bRAQKF1hTyOd2tVg8MlLlZ72qjYQ54GBtdMgb3FZzorq6Ubh437/IlBZx3LsYs85Hi/KSslGbktp
6rGDn1qWp6W/65DoAolSnzvYz1nMA3LJn/LbaQBLPZsNRYS48Kp4w8zJvv5sbYvr0pVZldqDGBeL
21BLrlunZ+jGos24WsU+3pAxR4XnMEveRXZO1i3Y7O97kj/VhP2BmqeXqw4XO2892Yrh5Q8h2eFn
KH5gepruIbsfaMxX5WQsD/B93SkIEK+5HBRFfpyU3GoVKDt6xlcQ5fcBheGDS2+SDhvnAvi9SvNY
F+jfvrX3xX3P5XkJopIkmW9GJ0TrP7C5Io3jzBwSTxztm/FEALB4EzQcC/pUcaB6//+jw37Sw1yq
dUrfzk9MILgChgZ7jro/1GYNHpnKkaIWcmOgHERjuBrHrKBCJnJc05VerPCepSLjHOXHltAwpv49
LOoYkICYEb/XHvlWAS1Rj+TiH9kozXzB6ApayLY+nhpzN8Rh85C6uuEq+x/UQhZPg/VfsMF2DNwN
QB1AswefQ5s8qY8yUiV1nHmFEp3zbeL8QP4LcKa6A87Eus9q3DDMZd8dWlW3MPX/T4BvW+l1U/XJ
NLQR/3arHdueK1/hpc6xSO/NOmMuRzkL80hYsqjiukmW2SidCUiBuaZ0LAkOVgfCNw0/YV+ecMCj
9imKu1kOqfgWwV8VvcIU2HMm9szqVgS/A17gpcd5pQdRZI+Ljd+4IuHmze2oO4VFq9+qzASS85hb
koTtMZ+Uyua0QoSR8leVnCOWBLTLH01HZhFqaNERJOBPhUS+A3PCWhMCGdrTJbgSbzOMapZVal0N
j5JrWKftXzRFHI5dLk+HYOrjHKHxHtJ67nUhyZokdLl+yb79T7muPgVXh9u6U/OaXys0YPY6nQq4
pb59LzHmN/mxqDMLNL1m+cEHXUGGFStUdukJmVDTN5c/OfdE7zM+2kJyQ8+SwFRCFCv6wmejsqoU
H9jbpS9m72vXzJkmG4mHH0KfoOf7K+S3Unre/sODhhMAU1vpnUu+2XrVDweKgB+key/9oVGs0PKY
7tkZlQiumnT+IA0FmwgG1r3GLwVDWNDEQCjZvLPNH34cLTMisqQJXkKL45x+/bKjvtsFqSoeRXtA
csRV5P75T1fA/Zp4XNamjaZgCNCIePG9Tlrdz8ClmUXru+GSqCr+6ngUL0RwUiT86y/dakewp8Bm
gpdEsHhsn4JpL7b+OryUUle07yn50uLqzYjjKekUiMy444eYWTO/U8COX3eomt19wAKFqjC5Q+tp
M1fG3rEcLkhp9Ww9HrFYre1ECfZ/DGzIrHykwLGilsR+uZdgFZk2wxscUNSDyl2RzZrTLpaqwRJj
OXt4wPps2lLwk/635AfQZuM3DC/iMNpBpO7Jk2PwwA2jtzxJ8HG+CD5MmzXJKwNMmYJPqxV6dRKS
6VMgFxrO22o0cOwkBoggvXOs+RkOp9BuG9L53qrOMo6bK1xezaDr87NwKwVoOtNfrNyyRcfJcNpD
jPxDUdu+NDRiiYAqSiw25Lg5k2vNMF4RiSdO6kE3OJEdGMdDl2fHlZB8zardysINJlP9D4qllK0O
bFy9F3T/Vg8BifzNLP+ok6HSbCjBqJXLbcz5s/24+8UNQQ/N9u/Dg/6YBVuBFpN093DwgkXTPYdJ
wQSszTABwRiObqvsrF5VXDlffBv5v192KDteNxIbStd2W8XO7uJjyHi7WQURTX4NV/1wKbJasnCi
RHmhPVQuOuPDoZRMEHq9wWIqUh6iIimwt+hpnYhDKaPBQdtYxEGEuzni7mNtLBXJLVu90P8/v8tn
AZbySS2y9or4uRc6DdzCcGw+IBk1nfM3DNRWvXM2EphenKTqhai9RfKN8qwFvT3TdH/Fqw8kYjlA
DO4joHDQD1QD8pY0s2k1Z8LnD9AVKNjBfGlHF4Tbbu0P/HzoYn8B+zlope4heRMIjp3/0zUZTrDA
gogwTyGNFpA3fwbDk5ql0J/5ejEJdtxGZ/08uQGzOZn4cIczu8kLhYEJCzFAn/6FQCfDl4K5JIVN
suaoNbQqaLmcxwzv9hPqlI3zFT/21X6HwUA1ZUwso7wxHGEPgpIgb3fzYJ1Uve0Q8Xl/H/xMuAJV
izmeXbTrkTqu87SsDwwzm+NGBktNEMIv/fRykq9LU9UAEwQQPV89sa5EyleucPM4iEOFe63IrQ/M
pjnpF0N3Y/LaX6lc/CHiQFA+fnQmfyNX7S7U4TzqaIPKw+DSn/vwll9UEIXF5NjBFjDxVRIQZqNd
To1+uukxCtXDqmQbXZDsYNwrnJtRMij6NOv09sHpecPV/eXZGTQ9AMMnvx8EMz8slkVFznBDBGcc
qZ4HuDkstWE68yvO7to02LW6VVkA0V1TuxnNrNzu/FXNUknIM0yezYBvpO6O5WM5nua3kz5tMkB3
qClpbhfIHyG923nK3VG1MSCoDjmDyKIR/DBclSh6qlaADerQKoUZyjtR8ZRk/1Wvq0rKvq3NpjZc
YFhl0lIayZ6DQVTCA0q+FP5LeFJhvRewwLLllTCE1HwHXRJE+D823GZTrWWwmNoC5ulpHehu5D2Z
xEhrMfQT9nxzvt2zFsxkCINUKq1b1VB6cDdIEiCTRUO504SLBp3BA6L1NwA3NpAwS6fKA6ub0LVv
sb62+o6V0vc8+/XxDvjRXYmoVsr39P2Ra6g5GnGZp4LwpkRfXr/YqEVRCdYJjmPPEtrD0+fxtZG/
IzhPHnPLIH+E0ANw0bncD5a4Tt4B99lOerVMG8xVcww8w+SsLPIa3mDMHZrBFAks5SZfw9aOdw/e
V6EwL8uI0jhdbs6mCSnYyiI5vBCtzIleP/iag2yllU7O/1iDfS3fyJO0ANqEEzcmYog2tlXgiRXT
5+bfdW/6B2ukSaYjp2Lt4IGjAs+akO9EVYjKY6m03Avss6l3wIG+EuoYFclPGpJuEV7jzQ5l+ZYf
Rjv01shXJMPpINe8mEoRXEjxAQyjBt3QVGdFAuilfeun9PasM3+T+lzB+PxiQRoySsLXsJDY5LCC
JPoLvWVyLjbHjgAFdwAd+Lq+QKI6bfkKkILbbEYPcinGq54swl0UGmTI7QlcVEjf+JcgIKRJomQi
kFV+EL2CAHi3ahAh2QHIR6xDIcd4rz78MihSt87kM1ZjUUd2z0IbqOo9HMgpK1EImr/K/Yu524wW
bBlhrVtgIqk4SCLVfcJsjotHmP+/H+MvBHv0Zq32agTRtA3oR0GKJfdwipbC+l9cYIwetqS7ws9L
+n/cNmCQ6EsfrKcfQqylItlk8JAamkMOxqI+KSblAfIynetZZz8DSGYd0fQPLd/cjXikkaa8fa/N
cc5CkWkntda3dUdujbKhZmyTPTddaI87cdxHbatagtcPz6CFGMXcB455+a7xYk5+MS+3LZx52vwq
GEC9zqc5GemwH+qmCIQNNJLcauZFrOI+dIyeBYpQMHKJb5klKm0C0itBAsee+L9C9PoRYMT/Z5wc
VLM0eoC67vNmbQ7OwZVuPufdBhvDGcG//8Cy1usek1wBgrir9pmearfui/xZbReEq6ZI89zM044x
yeWZCKLUxanTP97QdDPqJy16SV7MFvlX7avT8QHffxxkdQtXJreU8H26VZPugMvrZzozqmxp1+cL
Wcmuk6b6qUD9107EfyjwxCWX/6VKKUmtxRw8c1bsRKhiK4l0S++2VD4biIpOVsq/OWMMF3GXOyEd
H/sMCzFDVROYc0FVRTUn83uhgB9yvskYf272mDcDnCOW9ubSFdU3ilqqSWokNK6LnvS2C5I6QByH
QN/JqkXvWwkUGHmBQoqoiBk9ciHcDrlrfaYos/Hs777HsM0BUIDJdpt8cfrdUAwpBdZKa1Myb7iR
5b0glGME7cHY9UXKR6S1PuU9IhgijI7xPTyUp8u4WF1zZgGYI/ZIxZ2rQimWMFMj2ZLf2PfzL3JM
sOx8HE6rfPQk8UaO7Q66iCGsVUXQk08KtVmkCIfN356fPi+qd3r3rRa3eZus71zJb9glr+BTo261
+3aECDpma1wbINEbJ3UmJ1pV5r5SPUnAL83cVlw3ZV84y2TTzZ0gD3U41gDryJikRObhsFuTidMx
7MUiYw1a8fyzFKByBFOXzbhBPjrKElh46hZTmPAMGGmMy970PY2eKF9zm3u3PLkZZTqIsrPwsQ5t
xGxMgRt/0cCW0txK15b6BjBHaSielft32vC0KeEI9EmXqWWDt3ljvVJNudmV/xkwBmFMePYUCNiA
hqPjnlMWX5UFSFTgJesdTuqgJysOvtHGWxtizc7du1EUYXGXL0+SgI/nbo7AGD1FSG3GHAK9KmHv
ZHpw6LDiFquZ41gMqHuequxNcdERqRN2YQiiq9uQtnLB0CFYbdkd71KepaoO9RlUpGh3nPj9ZsFF
4aMKhzPvHpmqyzhLcGqYkO7w00EbKoNlXB2DgrAyXrO9utvOPmWoTy0+H1rLat65CHwE9Ain6wzF
r33tR4ijneWmcjuduy2bAfvjQqYpaazWB2rKyvu208agCXq/btHDsmppSiTRG7iqFYyrNQUa+xMH
f5nzgdoUJn0LXFHs7GVYIkInkRvYthDeAKeKpu99w2Sgro5i3WFFZ1ZU/VFFGa1Cfso00mnx7n3n
tW8MiKmynP27Nl9pJZOR5d+4C76UqEweBgQ1D+pH5dW+NzOrXXn2WirgJ4BYD6WR5rBD0Tcw4772
WJWnO2FVnF/MwT29tJlGIpzWUmczk8JsRXVT2zsrHVdV3Fr7jSZowxZfvVpkoC7J01AVeWoXm6O7
3EiPdBbaambB1AOipcrCDgohRgBuEr93vy+EuAzS+SWxWFGULOGL1szFDvNYp79vQjiMJex6hAQx
3dKDrADPkBTSbUg+FrQ4SnQD5IJL9ZJ6d3fG4MRHCz70YqwEmoPWTbKBG9iv+mGpA9QciAACYDQg
WYlMCq5soy0Om/8rz0JGu4+Gx74lKpnOIDLZkdvCCkTbGdWHi+0SeWniKoTUp5wLd0DYlF+Z6cNm
lznSgXj+K0Zg7b6nSIo77cq6HZv8EKyQV0zLeWFC9Wh/HR7mCXnyRl/oi6ArakHXVzdzMqSkkEpN
LtAM/4vrjqWNbLFG96ZYTrm0FAIlpikyRXQ1GYxKB9dZwAPd/ytvFaeuN0DLVTSK5FidlpdKaEw7
1Ozjcy1boeYkD8lAeN9oqkkBvMrY1PoYeHBF/eCE3e/lSt4ZkNYc6wfWnJkqwmxV/Ww2Odo4IOFg
vwdxap0Dd7dUDA120L3t2fPhZ9KPn8NrtCmxfKrn4ypnlNz3NZAlbv5NPqMJPOvNE3eongjJSCPA
zR+sbjrO1QQQNBDlKBtsSY/iXo+id8bhpn2xSEF29cJ+wo2iVrDsSkv+U9TqC7qpkuLCNcA2UHaZ
bIjezZOSRI13L2KwCmaSiQTTI9kKNC2ZHHT1vxj+UB22d6/xJP0LamvntcsLxAcx9ZjMw2y4+Td7
2M2G/bjURNC6hmkMNh1seCXmj0iHyinuUptXtS36BYWbDy+ZmSOfivmTzr3rv0Hhg3AAT5LWY5Qf
EKEmViQpjhYWsI+s3ymgzdY0OZvqqvpI+BNbcRC9b3r50M4zgSv1i91DkL/afmlw70XGlpgYkJoG
oWBymPAfiVsVy4gm4xJ0z6juYc6Vyn4sBHHbGWHegZPzQRXmd+xMaYKuyzyD46n1DjaidKQW+SuF
97QVWB+5dV6OVk9ZVNqNoPKu+9fz3NQOP8i2FhRa93Fq5RTQ6+UVxeuxyjUQ84s/irtX2SelqvpL
dyABpsk0KJttz0NuN/y5TSZiwYSOhNWjOhCbCZHZKh9kD8bXqW9I6cqXGsSdUoIkISfnQezLz6yn
/EbIhW84DTWsJO/gmR2e8uSmU78MMhU8Ttau7T8ry5EQiyNw6nfLiCFBlXbvJUMVRZnN+A9ucrqt
/ueIbi1RG8wFYlg5e+TU6VLs8TJMPdSpL67pJYVAjV0FUrgu8a8OXtfh+QDXcB0oiwED9VYNVY0z
53oRTJB5VyOUTP92gY85VCq2q8tDsadjtfiNK4KhUeDekqe7YQshYu7lIaz4Jrd49atJN9KBslDg
4apdwLdsSPsDrSYSYyIVdJICzIUeRwptvcyjL+tDzb/zLu+oeUB5iaCIEGFuoTgaowibE/MlHm6I
0JZQbIeZYnLQoJJKaDZUAozZ3eWZHqjCJU+GR2gh1fYOuFmX/v/Ha0zjxutQD5iSrT5mMoEKnWet
LP4C334NcY1EFilpQlQ5AMV0HL0CDvN7Zld/fbRmbo2bzqHuJeimHjFpuzOhlnb65MgUanmgYOs3
QECPPXa36OtregkKOARWOo1FDbRlzqhXfnZI0ElGhhSn7viwtxS0Kbzs6MwrA10K5DH0smE2uKCx
JzkUPMGGn1fP/bRfR4myIpKtoQ/n4o/Xlrp/ZIRGVvk49TudAPvnrEakPM9gjP0zT+2k78ifCWJb
RN/0a2fA2YJxGyCgvCla2pEb+6RXB/dy2rp9oeMp43OLBgHtziDv4tkDVkFeTkxBeeqH3/+y17hn
2Uz5DUY9O+ib/0+/7T856XVmc+Vpex4GoqsiQd2IQsSqaLfs/hxipgjRyMnjclCkHP8kbVgksI/j
S0n7bexRowEG2DnZOvCRfDKaWV0FPVwMx17HJmU/SWOu52y+JxKss8vs3DRBGxHBjCJCtQIuPfjW
GcZUhgUtfeE/eKKV4bvoD385Su8+AuW1DsWvmnvtbKFruoJhqf1bZgpg6Rx0B/qJq/Tdq9+Lnmac
0BxXog03EfWi4qZOTGokZZFRagfH1zWRn6J9nzDZGjlPiqEFexPxDlp16r09Gq/KeSXvIqtLrG8c
YPlgeXq3UU/qz0zDlybvW1ORD4t2vyos1m5q09tmRQxZX5HdcEQn1aLAmVpjZOqYra0thVbqGTz6
q72f/Q9DbNZB0uLniSXNlzdevSBbSQCwfHfYFs6ULRdW+vzsDZAX5klrD+cUA8sfRyCspeQs4Vwl
TqXieH0Xb7OkgWc823qOkjbdpVOxjYXo7u7QepDaqincd3pqoAi1+90ysw3wbKAGlAK69MTPxaWe
LYLKKEu3/T8dQrDAaUrkylYUYHf73wvxOo7VAf1oSNqjEKdaNoZUg+vPR+kcODeqD0QhOERnXB3L
2mPFi13G53A5kLUz0kHTA+FyyRkiZT8uROjbrjQaeEu9cZVKWb6oSMxIBjXjShxKnaZExjv8NY4L
wki0qvBTipnVJvQfqZeeR+9M4WS+9DFyvtqXdnWl45p1srZrUic5GqxvJQYKL6amM4BBA4U8178c
OT5Qj7xerS+uMMz2SHZcK4ZyWcI+b+SLLe/6+dWnaB6vzmBhJ5PeU50VbDIHOjZ5oBa4U0XPyovp
+h3tVtxQoIwSIGlaTzRBjeDXpTB0SHqyZVBGjyHO92tluOFk0kc9C9hWlgagK6PK4qMlrnkAnoeE
iCIfYEwF7gLuhErKCikMfmyxbjlwxFNXfnS/lZsrr5WWMqLcXFOtlSFJUDC5dWE5N8yuLUu5ZWLr
oaXTRoabpphZQi5oxSXjz45L5anrAxwrhrVf0jOOC9GLHfhfF20a+WMvt6UWnS5KvwLFCGZZ/Vnf
kz/BTYb+pTN6PvLD2V6sAEd0kOHXeQkSDgDEHPhrdf5OQYJCHl4WJEHeDT1HotHj6TQqIJv16LLE
Gklw/q5oK4dQvx8Yj3OeAQD0wEb/5HekkPtFk2aq6DY4tprKnp0lK5/++prWVoyaxA0a3yf9u12/
kjeIBdoteG2qTeO6iSTOoMApwpTVoe9A07K5QbYL/RbT6TNeGGQucOl7CNYULp7or8TiuVScIMaW
7JKOAz2fd+CQogYWbPa0H46fLGNwiPPFd5jodPhJuMqEPuuxd4weNJUw95pqEq+pOiniljPulkQy
BBQHcwYvKdS/Bz7ml4U5Ohv8//KWw7uQA1/HY2kW3lMBbDWBNvkliAllBQal/YwZ2N9Iry9q+s6A
W3vbL1YRhob0F7ICZPpuJ/uM79qgWQAwq7lUzr6Q/7zg4q0mtFZqzhrVGaBsQzBosCMIaeSbBZsa
rfJXPPnLFJm9jPdvl0qkKq+oda9NzUGE3Qbaheu2KU9qfyugZQOpcm032mkTPgxvxRDrAI10n/yL
mWd/B1zuLe2MhXT/ja1CUnWNo0f6KBThFAxnOKtTSfJzjfzBci1+Bcj3P+VMT8bSp4r+ArwRhmsu
Yuh2ve4gVggQQyX1QkJIADEQQcvhrLqBU5qow2M5+YFZzLfymBINBPKf8JqDbXBJbwUzXmcDTBuI
GxESqSXyj2BGAcdtjfa5ZMhTsf2Ap5SBbGO+h9X/ZCv6u6s0oUdWfp4K37S6kDAbWlSL+wIY0Olv
dqohufIpMquq69ONpFWPzD92M2x+n+Rlj3S05Gce2P239495/cpQl/hspCxwr3SrLdNhLI2U3xqg
7NtJhybu5DZTOkRUzyZJYYT+Tq4idJKqGT82cczl/B2asnc3XGN67Tjsw5HwKDscONwB8cQxsI0T
4VgcvfGq1G7v1LFaklqkaQY597NqbTsVOnnApktyCiZbJV7Uy8f1dN0mBOyrwev4YsStgb1+KuRE
zjh8EUNxZEw6oP8MMfzJ9V/J+wvPxcg8VsSFcm5UOWZcArs60hfFoDbkSczmi6iZq4clnwmWkHXM
KLMa6y8mpF/O4/CD4XgS6GI2OJmOuHat7HEjZRcLtILgDYX0RMKgbh+GogkZ5TGxIWJI3vrPkI9Z
8ZUkllW8ERohs2aI4e1bgBzGT7fbTOTJITNZoAbwmi2kfoztbtBjZvWi4OFlTHdJ+jsqJIe9c2SX
EQMFCCx0CB+FCrnKp8x1/cwj9elsEpq+YhCTdFiUcSOfJ73Akd2QXJeQdgCHIagw0bPThP1TYn3b
dZP18hYr1BffnCweJeFdNLhuC3lpd1NayDoEcTCtupTU70IqVcje1NhIWgvnXljjTSiawy0Ni5OA
27z0gLaC27bBHkwI2soXWUd/CbHUV/LjKCTVlGr7cY3vJ9quQbteHZ6iPCpJJkLmMRMivsivE8zr
JrqnNI3BGaIwJ+Qr6KRaC7DT5jDSnKHAljjqu6zZTz2gJiDZK2Skl4qkwDPJzCB99BIXYfthFW8w
jTL0L1lwnPpIkLyhWTwwYWcZJTMnqszoKSJ7FylMmw0bKDhlvqE1Uk9Ft2i3spBv87Sl0MiU36X0
ONqRFtqdI57S0fk1CzTtfg8u52lyNKVMeMRZ7tDZtgBwnO1rHaK6Gn/0I9nMVEfoIhq4T1ikOUNe
Oq0l49xCbAKC0kpn+QtEiWmAAAVQ3BbTvqE1J6i5xbQqkh3omU5A8kXoSNwIqRDzHN07PBZRdrjR
PghQAZTVycJ7I6jy3lTxnoK4p6TrqojjSPeb2MQvF8R/NWR0GD1jx720/o2jB5LiC9nR2gcCOLiR
4tzur94yrqqihBSkEod1RIk0Ps/a4mR50NgBbGa1CHA826i50JYev7O5J6ZUFHq2AueoVg4hIAWK
//Oy8b3/veBaihFw1hvykO4AOi1jWgJ/5x6cgIwRNHsnNJkXBv2iy8VETS0kfyDRyTpQMA4ciIII
1DhofRwXMjAgBtJMCMJRYasTbpnvqZpkhSKSfbeSeRXVxMCIdwQMRelaVyoAITyhigA6Uo7AEgv/
yJIoRojaDj0s6wZV3rqQGRaQElROsG8cANa/8JNOpyvttH1F0FzlRbDPyM06XWAckJDCi5dxHkfw
QdckGOneIbZajTOnXCLD9ltS+1RX3Z7pATorElVqAnWz2smHMBSHapC72/927gGIYkE+LijmIcdn
ea5jT905SNFg+b3UeKbv3FWwDh8tKbtbK0cGn2wsQNN6tsh4sGPkjzTfknUIrS513Ica2lGbDlZ3
zmOdN3WT3+Rdvhj9Nq96VsbkPM3JhcHO14FoZ6YkbPIJ95lJhHTEIOSpsrEjK20YmpG7gbC6c6C4
SwuxXPVBPboyo6A3CRUtzyeRxLpwhmkBa8BkRRAYGCfu7vVVXttuOz5uUf+87JILrsMqMjUGRU3N
QlhfgI7zGF6cQs9uG6vGGD5U6LHZfG04JHcSY3iFXD+uZVVUeOrjq/meIwg7+HrjmtV0yvMdzBd3
+RK16Cqr71nNeKvEdAhVtqopn0KGTkFiWsk4PdhJORrj0Cfmq97yPTmN4wVehZb3PnFPCa+WMZcB
GB/hRgzDy4S+6aEHBTYxRUqPxnvothC9emo0nCxZqFBptz8uVJV9COFZhC8c6TlFE7DXLabpMPwY
t32DJAJnLknj/1xKPSyz+m+pGUNe8JOi01vE4y80GHlAXGf9j8cK7maNgwUC13KlZtYATrfrjv5t
AP+5XHkz1QEm+OBqI4ji4MQ0FdRXu7waoetZ+zW0l7by0i4Gf3u6wWlce1VjtAbR6gnXQ6zsaCG/
qLgeiPCkif4Y9N6z7HrT887LvrIszt9n2YtZV0DicOukWU8fgzPSaXSrhtnt+lwfKJx7tWzaldpl
0Z351Pu/rq56nmkND9qAkAPf0YdT3dT7cYEAAUkMHuK/pO5hOki2/+hZKG0pLoghyD/JlX5nwKaK
Z69algRHI4UfOyJB4IFyiDnuQaDtljws9PQ3VAMjFc1CGj8aRTV6P7YAkQlQ3pOi50R5WsHGOdsm
r0tDMtPY5T/Q6XlAdfK+dmyj0TCZS6hEx51g11vfOktOWQBEdfrjYmZgG0MYfFIYYkxbzCiJHVKs
JroKuxu+iSg/bKGub08UKmeJjGIN5iFb4+tuICLkxojCUEVVbXCWsds2jnfOCOyv00LKOXTRZuTS
nTaZFWDcPFkjvmB8jEnlw9YWBRQUdG8nQ2btlNpqfkDqRXNuruuZUx4k12CasE4cp27CcAR2b0/N
jF6KicLH2yTq2PTLameLoPZvwq45Pbpnh52ICWEotAjOf/mNY92CHEUYPt1qCXCkRTprVSV7Hz9J
72aZHDQ1KrpGLrme70dYqzm84EUDw37xyZb8v9mX75d1PP1z5tEU6AECOIjAILzoBsS8ymT+tH88
CDvVdOfmOM8WQtJmFGZ8cyK3G42UyhqiiS3YQzRbh0F+PAe3mfcNTmPInz6ZquVZMRAIHLl5pOoz
tfESw955ZZ7+8704A++plBPnOSfvY2om/JT+rPz3dPlgRlltfAuIfXbm+zHAyWFjoETU3RZ3fOpA
z49Lx4kamI6ocqKeTEu6ZF7R20zC2jGws/4MJi2dAt8SjhzwofHfjlNosWA1+i5yHc+U07NGiSBo
jXW0K+cP1McR0JeXcIHHCxxkYK+h+yMRWjml6FXcnazx6W2Kqs2Z+2K7Dae6ePU2sZ0JaoZplDGI
T5RTDW+59UvxL/0BfTIsHbrNmdgtPqmwxE4nkwTd1vM1EDOCxQz8Z3NVSDJc3FRlgxqjXxclLubH
OgJh71P3CUqhqdnPRk86GJ5dVNDiJ3Nxy9eSaLjuhXHAWrc98ASGzkQaYu+Vi6dUwnBLiXUF0tkl
NIn6icWSoy3VTVX/G4u9qQuMSGoBGI+zf31siJHuMG0BKlVgqGUiOJ3cqsk2/9o94ItqFmjw/zfk
VxrrVBa3Tc/RF0UBp2ldxdKnn5ELdgLPDR3s7JLwiZCyBfIyT4X9eKCEmaSJyAhOga40k2HUngN8
Y0azXmwemciubKtJX0WJZ8Id9tBZFHSn8go4byI0YQXkRsP0ARkW0npP5PlVEKyHaaFldAu2g5i0
8otsI1+PKTXtiCm8mEa5o8cLZUYAdjnSXVgtCS33azqmdS88Entii+0SdbCPZiX81PIXw/XcTxNA
g+GTvIH8/xX5YuW4oYyHey2aZFc7A1WqdE4UECB0cAZqHvwpEvdJbT1avDfA1n95+PNe9mz32QkF
Qrs4yh0eV27PzMOPwkQ4AuDMAywk1R9XPNQaCUju7o2iwAtPIsmaIo88T1DQKWya8+rCVXtHKwZb
TmXEMKCoOCd63xOWbiWpDvn5c5kVOFHvfB+Lt7d/ZHrE16zJ55nUmIIIhtYTEmxm6c5+BiDXIyMo
9Vg0vWEsVKr+7kX0SexQTLV5h7qmjZS4O9hf/UvoYRFmGaUBJ7K1MaLRI0UhCTLfZEbTKQuF/+Fd
gfFwQPfRdkBcibl4/wyzvIMejG4ET2Ph9IATBJZrmv1E7U/3SVmgUwrfCwHsxuw+S2Tq0GoD7Xn8
zyAz+eO31UaFDB4d1os5JvjCyO5ZnFSnw+Sj4ZsoxBr6EOaDb6QwGYkarNKBcr+MEHNdsVUmRF9h
zCs4qno/aeUKOJKvU/TcM4tTnqqVafv0uq9RJKd6ZIDdo+BEi6SJmDMHekMfzAyk/nQ0Y8Ng+qkA
LBO00UixCn96p7zsYgonaw4OSg6CqIV6x2kvkA6K/5f8HK1kZrLwJQd162hc5gYZhRX57cfBT/Gq
ohg4ioJiqNrzIY7XeLoncVLLXjqUrVoPTGEoL8j1irTKc/flAeBQCgxm0Hokq4aHNA0cexLqsYDT
uCP1720d4l01gjiab9l48YCD9PIIfeWJ9GebtXRktG2KoCpltdKtzGdTBA9xwXArEv2/0P024eyl
H54B79RZ9JcPX0cT9cHqB0GQ8FZ61TVGyYt8nHDsMMHXjMDiCbQUptxBvoa9Nj1mC4JF5HqVMX7/
2215/zEXJv2KtWmpqY4bdxXWZmSW+h3HMrmYmmXwB/yVPACk4hkZQZCIHhevn13eipm4/XiESyQt
qrTAEs59K7LjNN2qKYXxHRziyT4A9Oj9S3cF3PQOUFODIgbNcsuYi7lpMSjGrv1Z/irroKYYp3Ch
efVTNL36SE13mqRZD8kiksqpWgMNVQoXSRRQo/rR8PR2U8nbmpiJ1A9ovG7tCdWh2F3sTqZIciEN
B3Ge17MbAxfZYYOg+XZr0MPFGM6J3/vWiygkqHy1HGHeCbqeOn+9noAl5ePldEjj150kMiu1xB2s
Qd4MZClBQ7s8vPgoamc/jem5DPHI7KGIJ/VslCfXGm6mSzOMnaGfBJKNvempVGYMnrmIyNPVpJl8
rvP+Iq1KYfabGHK5rT7OzdpZDQ6Ta+k/o3hSfpZuKVWvqYSn4EsEwLMhiqbauuBnxUiWa/pswkjY
WHoU9hcDZAHfwd9lNvUBi0hsDOxVVghL6oXvcmC50T0p8RadcdkrFNy0M1vIladPWM5t3SpxLOr+
NFYrSkdh94anO9907cieCTvE5Y3QDSArOEK2nDuWuat8t5I5tdYQT5P78xya1drqY5nNlIa3qMt8
Y/FMmSRu7Excthqk0DBMkHGWPvcVEqiDoPjL50DemKHMnHiX07OWl1oI0aEYKTnaNHxdHJMyt7NJ
PrVckqMd3yUkI5/OiC7MTCah6FaX9FOq/J47x9YfmdjqarKT7xA4yJzwZ4CoQpJQ362huuLwlYPm
QQEKRfKU6NoxiBVMypVuyQo+c1QPVvdU5uPErOfJOiIzLLgnj8ggHAoPxO0XNYf/vxWlINKMqTwA
oVQVlx62GvoaYjAm8D+hUov7aAAh7KwrEmrdmaJrGzvVzo4bqHsy+KYB0040E8wS82nt5WrpMv4e
LuRVy7J3MULNc83HU8XCZBVicf2dmJUGhhFaP3wMZGjv+vBnNGtCt3aLgJGLv+UldZRVC2dibcRU
PA7z8gg8f5ax9DX4GomKohzsC3DkHumEiR4FJFv5arFUbE5BBvib2ug5odJ1BJrJPjI84P0mPku3
3dAeqsWfDH4BKCuwurXx/jtDR6vOpv3emtZRJUnAguYXNlvHdr+xDXxXK2Wa8oxKLT/mRMzSaPvf
FAAH96PFskQTh4sPLiOHFeGLZ0CYDz6AyD4AeQqdwMYvTL8fX+4+8TWfQ0Tk3KzF7+GLYbjrr7ZU
RCFVZSVAMvqrN+GiNk/19zz+sK3ECVKa/AVWjavDBVfCRHsENyEOqOKYQdmWvrvTPeUskJ/VZXiQ
J/9oo1IBwCOzU/Taz6n2gMxBo/YfGAfHKIsRia3Fd4LDvMk8TSdwA7crWMuW+ICWqmCh3lRTy7ys
Qi+qwGxKaFzF8Tu8j+gJ1e5XioYMJBVyP0xFLZjYrtSyZj2o8WFU1FgULhwjvRUJqsTKBBIX2FCX
mi8rHqHJqX1zMz5VbUStQLgMpNnqcjmcG03twfETuJ4xcQ+2xfZlKRtx6L9OS1x9R6KQsf7c0P6o
HfTZHAFfsvghfO66wQKsRHcOPrHpm5D2z3H+icN6zWqvOHDyKPD74UtqSao/jIw+xiRJFWS28hTH
3f6Zf9LxuUbehC46E1xKK8aOxj6lglNi+s1AOn6h5/Nsz8dZ2483Lz+qLP12DbX9t/jhpBEaLzHo
GX8WxYlF2WVsJgmjnLMe9RvCO0uu8dmWcYFyku6AB69Bn39Fve/SoydB9gJyQ0GLA6g+bINoqbo1
M3wmGF0V3c1WJdYcx1CpRuIJ0hEMWkeVtmysohOBynjck1u/4vca3CXOhRK3klqYvLpNCpLA2goi
tUrJ2X82GjsRgJEgRbOgzlCQedXhkDpBlSz1KgYpqlLWc0zuYyrTvEXO3k1fHs67a7GVTr+yARr2
2I886PCA9SK5E1Fb9lrtN2EpymQ8hi79sKY/OjVzrpjt2Yk9c6a6RD+y2ZynujK2IDjU0aLO5pUc
AstqTTL9DLWh2bQHwQL+YC48N2XXJYv5j6fIleV0miAPevHP01iu/L/OcKYgJEXesD6CPcxLXb+p
+O3T+wE2Uek8++L6IQoLEkB4YYxyYG+OWDOmrqZMXE/1xDs/7WeeStf5NdxPBH5zW2iuQBPhbU+s
NEIXD+UEg9IBKIQyS+9O3eRKeDHGaCGmT2SMCzj+k2oxJ7/0BjAb1jBa9hkzJzqZ5ygEi+CVY8E2
7QsWXrYP07Ens8PHr218vQU/XoYRXY2I+RQ86/WjyBLl4Wdk/yYq0PGbKXkY1FvmduIj3vX3JrQu
l2sfEqPAX2TyC9zgwsiIJSvfeA0KZw00TyG1TdG9jpPcWsXiJmF5cx+7OpyG0rwO/+FSxEtPkVTu
ffziO52cVQg+Xmh6Hq/sfk8YhC+ZriINVx06TceNsLiLYHUE5bx4Lg0C5nNkNio03q9vQSqkUkg8
R+ZbU5Es9fM7aHI4sTIQ3DuFawSo+KNsFjqw+LjKsad5BRN3Fkr4MG8gm/aPj4Cced/nMLZbfW83
foz96dlGsARgvsPMbrL/a04aC+p5zcXbklx0iKviyZ59xCTRsuFFr27pLEPXFuTKwgE0LNsFTTKw
pVLYmGDymWxvb35OL2AYA16KUMvVWFbKsjfCsBLQ8izZrurB2cM3CPwe1/ItQsIzm4UwBoTCseXz
0mZI2bws0cgJuV+Ng+Oxu69oTgqptbsA+a4d3XEn2+f5re+qZPkc3JFVg9XAWi4qiPm2bhkizmt5
B2KrDTAKV3JL4u5lgWf1FXb3J1XzJAZY7OQxIeWEx1A5TAf/J7JnLzYURGkb5GtQML8r5sPZPE2M
POSzmgaH8HgLFuqskhf6IcGPabnS8bdwpI/47oUaoo7gCkX0tQ59AxEO6r0HtV5T9oDjUaawmKkz
DANMWYPE6xtQwKvMbHmb60G9gJA+NTFwFORxX6n6BdANAqbbwEf96KORO6s8SbBAqSoRk5f3hiD7
rEd01c8PF0h/lcES8hdd3C3r0W91bLeaeON54Wl0OGlYCaPEYY8OSTJJmgOIJhMtkswI3u0rc+Bc
D5O8ZtJYuPIljtSEhGEEeLdp+qOIKzOUhwU0zsbFFpdFuatkLrINa+prlXc65gV4MUA3b0rLuhGx
Nwj7We9dJqIxZYskXTtPbs8i+13xzYSDBkeRrnXk7tL177suL/ZKUXooEICRD1NDt6S1p7i4r104
0xW/J1zmHoCtDcyINwsQRSRreYGWJQhcFKwDvZIFaIJ7ObQGor54pLcaMtMSlyut3lAWLU1qdyBT
iOMggPTabopRDHY4AYCMgslSNlNULj55cIa2LGxWq7glLFbT2uLaeqVKCwjbauw8rGCN3ouBi2kP
pxp2Jy6VCxKRwYvF/4vdmdjUM9wq6o03UavdwclH8qY1TAmGre1MJw8Jfl2gHaxHSCJ/smaOpAnt
/7M6RIcDa4iBlAPB8CEAwJIQGul1HJoPab3R/X+WPLs36Oy5n8g+/Lw7W4v5fdouQlg31yBFPcqF
07UN4lFEHBmD67zwPp2C7WUbXoKhJBcTct5yZLpniRxsLHXPLps4ZfdVKfcqv5a7Jh5+ME69iTjA
ElYlVgw/XUzPO69eHZwv4+zlXLA8dk44HfyrzxzS+tF91GfNXUjNtkUeyEtSYEKU+DQiBQTJ8Hkq
J5//4/PsuVR2/5oGNRiTyA1V8+DrccFdzFPsPfp0iGo6r4iwdE8nh+jW3IXnGbp6CziFfLO58GTJ
AjG+9HNVni+ZLPTcgRU2DyKMNPZ+4yeG8bG4WTld/lB7mm6S3vKvVWX+mChZNi2pBK1Y/95/yi+r
GZh76GN74hZyDairL0NtVDMnnu1s5D4g5nP8ijyOrfFKuOYERSZkcziyr+dgxQ0m/JtGysH++uX3
ivL8co+2Dgu3pjm23mO9L0BBBskRzuItOcEQEBPjFWL91Tdq/DTZ4qDVpb/GV+5Kn02GzF2q5ylP
O3f27RSoVu8NVsF7KO4TOO1odOvAEAKG2VHRPYfueseoa511064mH1smqh1mo85JGqfaWqIacqHl
HMDWTR0MEIzgYQgEFcZ1UEChIHWpMrLmJCG/5UgIEMmtjDa03yyY0fvLqCwqFxbp14s3YoWnRFV6
pDGhidjVvKpReVRLE+oGrOdI4PjX5aefgr1o/kbj7uXKC91rtIx5zyy8fKEyRQFBI6dGoYzko3pP
Eq1RT+epUE+tYBX7fDoqvqfJ7T53Z+kWwOdOSj4D3WoKEn34nd9WA3DRKTuRMaNiHSFvI6o7fe7D
FITPhawA1ZJ+SuAhdiPFaDMVoIRRSK9zQAx607vt3wzY6fmC6WvLnBeVcKZcTfSuJix19zgvGwfp
nyisXlGGbknX7Q478NlZHQBqcLVG+ukS1EFbJGK3xHFjQkouTFmhoDX5vWVdhUlYAKIOmWFARdBG
/s7pdd0B2RY5N3CEI9CbdCfUzPg46TACu17qqZMVYQ5IBQjBt4l9o6RVzH0d0rq5shq2GewwmXFY
d/Tv/aZ11srUJRmMBP6MKyLkPOj0yyo4zoykEQYj5lQ/Wsfnsc7BDZ1NSPONnmgV/ZpfiGhNZe4D
t28SPAYfr1q5d1/wyvEfnZNvXhlHCUCgdy+XiCg4xKUKxifuMYzE+tmgRBweIhUclN3DRfQydwtd
1ZjKXM/ojAggLbSgYW+IdR/s4PU8ZK0Ct91NYq2vwrT5GE/Qehvg/kpCuPVBwKfcTwi1Ro9tlmLA
AUbB+uLF7tx6Mx1IyyakyryzvDD9FZJUI6p8+Ezs2eLhysmvsTPh9OQ0NYvborkGzjYerloVgcgX
HLJMhDtiCkdiMH5wVrpJfhRNIqLRIFX5DVoeA8aKiejCvQO18J/EoJQwDX5kndHs/0WYgUt4FP8F
xlE3SWcgdYAEKtQ4uVaPlel2xCZErO4q8N3dt4d27SPUktOZpfyut3Vp0I8gdUkMiP/i4sGcbV37
PH5XshgTNQsASXYKO2sGEEnDOWAbAXOhjbtGfTZlirV5CW71eJzHz6K0Sx8ZQLzAgEGgPi/0pwLf
hcEQ1G/UHYaHQ58e+nZaFRlqLJswRqGyugdQnRC8TePEgScbOBYieBgc/43c89gRsSyEoKXI/3u5
zYn8vc3YQ7k2wEvhSBD4mkiQxjnxvwFHyQfpd4bQ/wcrE4gnN340iZHmgrTgXgCTZBkQTTWZ8KNK
0mrHDEka4XsG91rzFPMqGz4Vkmv0zApG3cNRsswJLM9P56E4uiCW9/N0F4sIZ2tm+avJACLtMOMc
iRyCb8HODvChWOO8qoRBAAo+xwp3M6k5p3y56oIGWhkJGgmYYVZ0b53KChUGiThKoeCUdtv7DjIi
h2BtDgtEUgPlFvuOrmGuKUPFXG2oDRHsv5Gv5ZGi+SQUQtmwghkqdyWc4MfgRI8EF9NJrxxmW6UP
+TIDLBufujSKmMwuMB3eo1ISkw0mocvl+lC7hltFkd1sJB75n2yo7DUhqXlLBXB40z2OPKRi7dyh
7eB1raoYDpUucBmWld3Wz/J6b3DO0iUZ+UPc8wzydzXY2ei2xQMyTUDaRPQdZ+w40dBrFSRmrmfO
hFmoLs3HZwowrW2z1hJiVkCgSd4w4TuZs095FBfvu1Mm/gdayydWXqOehynDFlWW3M0tSBalCWH9
+iZPAS96XndIRl7/7SXMYYG7hdhB44VAI9QRVYxFciZTkZ1IwR/+9D6eM8BiVgHKN0dKDGsivVBQ
K4PYy0DIXRSLHy6q+Vs/2QqsShpxadnlkxiq/6yKI/mUhRj5WQOubXdWGMWlst1oZiwX2yyC0yJf
TKcUzjxvURxQ9PFbr4Gu/VkqrgqRYamGNNBIjJPL0wOYWe/GOyqLxOu44XqnJh79KIxvP485uXTe
Hq+D8M0IeIwOBgXUieDAosHdWnZNioMANkROSbzqxL1kuh3+GzdG/DtS5loIS05lc8lho+ni33Po
8/SlF1E+Ao+GqA7t4fOk7dqdJQInJf9sQzFHM1yObn24dVRu3z8Lm0m05rsuhljo1wJCOP+yuRlE
y7oaYuS4eam8m6pFQKrhwKCHU9YlM1nkScFCkCBb1LA2UTuEeIzu4i4ltlX/gT9Y4iZZNj5HCCFR
02wiU2GpkMqFGfdqRDVnibOfKK8vMCkWHzry6zoGQoU1anjdk9arS4T+r5j8Z/HN2Kxa8fIziCIX
14RTakkRIRE+oQLb1NjurORn2RACszaiK17IXa3KR+oDJZRRg1rNLpn92hhcFbUep86ZYWZBHwNq
Q57BfIJskCnaD4qRi733dgUjHqvBO9lEgkoHF+sRXap0hy0x3BlXP6eLCZ7+ZX4B2QsDX7iXCxtr
VzultQLNTSvo7lvfwoF0lM5IhOKYUvKbIHt4m4XRTGAoAy72VfZ5qprU/iZB4wbfDn2W7C1mqvcN
2W5u+omiv59K3FaxJ3uKKTw1E+YZp270i92vRoi15JmNoxq+sBuO3Rb4/fBUlY58VVoR+fgMDe/A
X1JXt2334uYbDXGeDjs5XW1iTq1Ca4l2KG9UAxTuwyFObFRCU0Fxwtg5XV1PwgtdjeY8tEkMtowB
3gQwIrIDrwkfA7yj+asogkL3+x8/VQOLxrQO+9LAC34JOYLG13VG9n9oNf4G/27mC1ykUXaizW4q
aauL2tSuiGXIZfXQpfuEYvZZPJfhNasFxAYDGg5ReffKXrQxr6GciKeeui1MsocKVv+kq9wH3/Pt
F31DZUp5XVyUpQpby8IJdsM/JSl5dX2JpFC6Wk/WUgnaSM0tvA2OiEz124gFVF4deWxlNH1lRzhn
kmebvlI6InPcWy1tKeR2OjsglelSSqwvIKF0Opd1hwTJ4soIou5LpJApN8uLnTfzPhVD9LkQEK+L
S7Nvi24uDr7dHbt0tInqpx6A10tOoZdQ3qk82dfPtjd2+d+iaKIb/e/2YqgOENlmSvsVOniJiZTy
2x9kvcSq2VXMAHv9NrIyuu6wVsw9YqDtJzmU1jw55/g6nE7ll/dIbKHvAw7xgdl9LDj06sxYZvCD
G/lEfvq7aJP8WPb+jwBNfrzrDuR0/ljcxba2GrbqRz9kVxGWuRA2q+snVwKnkroazupZtsASmI9r
pUwC9JtAMO2NSe6wLtNpEwPTb6OPO2jQK58QlBhMHSgYhLRNrua8fAsv2zISEkLreIT5OystOlNT
RFbclRKZjEJ3qMqNSqXXHrQ4chOyPYmoTsZSmMvNEYSQtz1zip4MFsFDUwybf9s0DrL8J/OCVbkF
wBlOgDjJuidDt24f7U3sxwusjytOWG9GccPJp35zIqXpcsGTASwgQD19zVxA7i2VjPusZUZnCrTx
f+kXWH9I8Oo63tbk2yFxcnhoiRdJQroU8qDDUDzMHg/zFXlzL+b0P0wDL7JBD8hbjU5kGc8hyqON
UKpSpV9zn2S3X9xpwAr1jZX3GWhGQgpz61A9KsjTI14q5aDa3MjJxczPY6kPa0eb5znLS44pOS05
BqNe7MFsgD17JBBO9l4ZWrA69itBdIwYpddpxdHQ3pMjuoOH18NaWghFGZymHL0GhjnnXv72qcQm
IcmgzxWNF1r9JMrGy7YqkvnDjFiWcG40WCqon6Fk1Ope9p5hi58nfiBy1b8MgUdGrgmbtjyZOXCP
zugqYdDSyJwJahQ6i6F4cJioDRKUsnrIXOltXzcr6lEmmCveKC+lrNxIiDvCIrtaBsfnvzR45nSx
N+SH0EpPOrRr2Dxmiwun9eY1Goc7TA780Dj++02AlHlIst7GHU5CUWkSXKB7tqOS4StlVdIpayjg
xKtfblg0DojIwi3OxesSEhewQgOSruxH9H/aMp4CUVlTnFHv19/LYLXBNpzV6Dqq0XmKzUekmPsA
siovYzZGQX1xQJ7ifr7cTQjeURr4m4+Vj7XH6G/SkTNEOwBVFit6Dx7kjVbey+3TsPc+t+cyEsQX
0yRGD7NIzRheeShw5cFtd+etuWIxc1QhBgUkQ/POMWa8C9qRjUjMrLX8Yw7ghcO/y8XHGQWFXp0L
mBsBHn9GiPkuZY91nDd3tb9tQiyyMO+VLhv2pJ/3pZhME8EASHUkQi1O6CenfAO3tkb8F4sYlyA4
sdB+f2z49AQb4M+1aEPtwsTx+HPJb693gKXbaAShvJK8lh/kKbieo7ViRl7Gt9WCqfYUd3HSptdy
S04CC7s4Pvw3cThQz71UbS1csHQcK5fgUVo30Bshm88+v7X5y5DeUIYYA/rE2HOs7xKP+NvmBPFK
rET9ffDon2zPM15mSIi85Jia9YOyq8zxPtM3Bp+k1blbYkEKxJwjgNL/wmjMlnTxyAdZNohPeBZY
WEA7dne8EDZKrJFtmnisU0UhAAj7vD4yzAW3IEi7Kyt7wO6m7lx1wQypub1uA8iqwJQDpt2pstWH
rsprtqyERlxr1vB90d+61R3o6V9Xa7dbGLAoWT5QgUWjnEr6kbJlOUh7H+7wyBoRRgAcIdkU8cI2
8mKF0xpUc09hg2dnoBAbvSqK8mXca3Rg80+C2GpN3Ukg9h5iz79wN+wQRfNdmx4RZ7VMlcMbNRPB
qahZLbNMEVNp1rnI0rp0zzJ89wdz3t0Bu0YnPQO7niIyuuRc+l5zqDip84xgV1TRQxOU7EHq9sfZ
fuDKSMz+mZpYZmRrW2EJqAOy+vs19Ngf+oTyIUF5LSHp5L1xSURjp1iYHVgIgFXjjk/xSg9HLxku
mF5CDlrBJc22xFVpJxwoMjLKHUOks0ZblGB9lp9FAhXGbjRGaiHpmEB+7TC0TjweJTE00xJXDihW
mapFCqZ0xm4UAb6VPO2uBMKujM6f3npVpRAqVoN4JaC+o+m0wIvwXTZIoNbPVkyHEPEKwvuAGSm7
ren4basxcWmI0G9UscJs80VwlFTEvDay6SX1xSM9oUAzEx/iFWjIKbmDWiDW2RTjXI2kC8SmJZQt
uZ99QEULTaqTy3nzcc4LKoNmg7YRBwm84hlINWaw351UsjMzvfaRmhmpW23TEPx3e7LiI9hSHKO5
l7EB3HHlEeTH7D9TOvt+RXpMw68jfzneecPbgw2cmElVqTc/OwDOaOMY/3cstdwtezfhwmI0ryyc
FzUb4eYXt4wFEKzvB2lA/W+FPbi0cW4WxrJsFaoWRBux71lje+Qvc22o3pWfBdlaKIBUMejT11wo
9pM5f0EvibjEmhwVJp50HgNbXNXyN+zzzgyJmkeAUX9rl0snGY9tdXAsue/uBj9xTZRkkZ4Lbk7d
JNJlUANpaatVenSV4zzXWFmgzTYKPKYV/9F4fFbuQuExFlnfSCXi3Wacp3lhPxpeAAAoKth2jFhu
rmqXPYojXpYHx9KtjwSK/VzZFUl1w3PfffdZnWQ9vr3JCvmeNMk3IlFE1h2QbuF+OQLCuCtohVXw
1Pd18bEpihth3bwWFxKXmQQzXMQ3+sKzPzpM6O51o1hooEuQpKhyNdRv8FPOAeLmikzNvEIrvpWH
255CEigTuPo+CDxeOPfdg0kWetdRv3BdcCX1AzuDzHDP3H0SKw33I7GlLmeOsZK7iL9Xl9U664le
2bSsrUC9ynj6tOSmo61NLek+ZffKFO3Grd1edGpvm6bBkwnDNcivDU6iCupObRwvMVZ7naBBfgD6
pGAcIfIBOcmKYqHV/OCfGEvU5C+lJ7A0ElIzEIsBXqdvpiauZm2hb+XczoU/zP1DGjccIRRc+DcP
NFbQvuhe0thKPeZIo3SBIqje8Kd6v3DDpIp5JW3YUe6oW6s/oKCdB/kMXQnvU+fJFW9Su/RmhMOe
GDcu4NdnEXyAfLDIPWp54lXxWAxbE2TYg7dG6lbilGTiJFYcVgUHBEFqKHohHVzT5gOIr7yE1cmv
uEWSohmD8kz4/iOROmE1qNU3jHqJOaEcHfJxaOK2OG+Du8yxhhwv4i8heYxhULFrnsrPTuhDRWCx
gnSgAXTMrjSAwie3UAm6le5q1vi/+DcomdqQmwaiKAfs6afy8Qosp1Iov1vuTr4j28wHDe18GB69
pz6kCuMkaYpDG7GBTTg23szXOOIkMZVgT4FLu9Fuh2sx08ncW+xTaCZJivr4yHp/ZegxVMWpWOWZ
MB38Wtcrhe3hr6dRIQuPUZcaYx4fQ+cmKdH1id9GhQykUmzlXOqgbdT+sOGdQJyUu7xrLYuM0eRt
gnVpFUNEY3V0vyJirCdeZQcEvkafsIgI+sZtxgF1GViRJfWu/yNMg+3fRVxADGCXDhP+ylGKjkkf
veP8Mciv6PKb1fKq3UO3ylFDvk84HuvZvUB53kKlDOX7XQn+M8QOlhAoM3jUB5Q7sdeTGKXdC3+4
yoZ0UfdoBKg6Rmiy3fP7KoEfYJ4wgsP8JmsrT/D6Tdwid3sveks15oXEWHmB/HRzEboi0klG1tdK
8+zdp69Z1DMt0va8eH3BOG6BzGL/2TCTmM+xIg6xSU8FjGfK+hOCcwfk4Sb4orEKr/63Ka/WvdPB
FlntpQs24tWC8mcYBXdpx/0vDINOHItUd0FxeQ4i9H4mvrki8l1tRz8Drx5ymu7RbLNAoYPQvyje
dWimKhIXAtEh2BrJKAYnH49I6rDxbrYcXQ0GgOk1Lt1A1923Zdx1q9iDeU3IRM8s8eCH+Ai3JVXW
diCPrsKKFDcpEU1D2E2MVuEVBssRon4yuK1oIhK2oxD9V0nyddIVyaVWEyx9lyTvR2FFDPBc6dC2
0Alqhx5zBl7hOLpmFnyF9fGksJj1rJyabkdV1Gz3XKtVgnik4QQT9XAXZCJ3ULUv38krUABgLf+u
mGnzgNnSlzP27K/Nqxu/P0Zt7AzIvcxcOhuZc6FFABhE56bqVEJaEgZsdnCGej5z7DJ/qp1xAAVm
X8OrJybFaFcHATw/Pzo9sPqZsNJdgN8lhhtG4bHTQ6UCnBQ2K4GFKWZQ35wrH6i5LGapfRRe/E2I
5quf4lv3zVS8GTfm97nmrFtk+ZveiSoRPeqXSluYrweOLXG7j/wNsIipSYKPq0DalMR0PLIxY1hQ
F3O6PMU1yl1ul1zZSgqxZolFBy1xT6eLIIjJ2OVunhMdIJLYB/mg8wHVoBHFa+PrSPi0YA/pUR4+
pqyGLCYi06V5qvlgKfMW5q2YkzD5H6dYDdMQzaLbNNjyUI2ttYz+/rsx4VJr0Z84gPuygQWBHY/u
HVr97LFA43cI+EOGvuKZXfi/xTlWgSVIrNE1psOr22nhhhK7vD/cdVc+PlmuXb3J3nPz575BstHo
BJyDCf2EfQL+prxmiqZ5hqw4fOG1uPsEWtKMVKFDsghL7Fu2EC2kvaWWcFFOCcz0cfPKpuGPCUQf
/JO/q0U2mJmADeF1tIE+fd1KNtl6uk8MjP4qR11ysxkwnhdVgV3neoOPPGiu1P1EfNfHGoIANd+j
nqQwKSvko5TMKwIQfJeO2nigOAv5Dc7/TfRkM7TcQ73pnH1aJn1hf4xiHT4kXroW1OH979KytMzF
OgIdpstERqYrwGF+By+yx2K2nij9+D0pP7G0xFnUeI3jjhKBi8/fNrWmrYzxkWhuAbxKI0gYzPLw
VacTjFTO+Y7cLf6zXWx5bBQ0UqE3IUZcUIWbd5gvE8Qx8EtF4bG80K8aZ2SonFCW0JT10wPTmazQ
xGY7HbBC7lS9vH0MdokfgyPb0RJxlUX+2yuALfDbYXgsMzSE35i0xAEUvhS6TJRRgnTP7FYIHNby
oGsZaGfqNCOuUo2VUD3Aw8N6BaRk8vucGsV/51EikMHll2IbW6CO3XMQoirYJahtCKdbhcZeLSbj
63ERSku/n9Gxm2/67kvf10DWIyvU9hOELqYhWaaecZhaaQOVEpmFqLLrVK7zujtCEKu+O0vsFAxt
ONpmS2iMDylKgCeSjG9l4Qa7EYjaTe8srLfwN56IJxJ17Wc7JY4peSsD9Hm9FWatd23hx1i8Piig
ld+O5ENHeA7jJ62mPXK7AqPzJtCKaTirNl4OZoPxyR+DvvBAPnq6H1xMMI9Ojl8kqGwUvJX6ow1G
Q7/QTeWXllGVztKoJ+3Uj2qm2PP5cWG8MA3amJ6ZCOTeks/MHHjjDNjLB8a1TssrUk8C7aGDlArq
wLe+Mz8WmnqfvIITIzjwNw8pZxaEi8p79sKNgiQkmMtfNAdopGZ8FkJxfMZC5X18zKSgl/wAJ6OI
h9ltEGlMQU7ltlQoyHR3bGGXFhPSbBN9kdfmmxCJoYv1eHEk34CNxYhye0lIKYIPx35pkJPMM0p6
etA5SMoogAG2bDsgUBlan0clk00diTT/Qio3Ya1o95ZJ9CiyGHTbK8KtD988lJ59e1XkU87hQrqf
7zYuIEr1fwUrobPzByQEYdyoAOxjcVhTsD69qz762XLxYxyUOfJqsEZtCYiuc/k0O4iGiXNT6oRm
eCgLD2K8Gvk5wQCETOeelErsnYzvrlNOcXV2GBXYkreIxQmURo0IOdQ0gZ5TmiI06b04ybNog9x4
3oQX0Y1Y7ivEYq0kRY2YQ0dBAThjHAEWuwdp/Ql7jXD58xow2V9maTb0rTnDR0wF9XcO26TxJlvH
wvopcQvVSj+mOI4b+Coe46Pu9vCTM5i6f3PSRXNeg1DFg2fPf11sBW2sk/giPuOZ3tzm+uiW+RJl
VkRGCXjqBL/6t/nLOkvFBS1W/uc9D00NCOsVlLJ5rot531+Ir2WgYna3D3o2r2Zbazt2XsCg+PoI
2CAW/vbVr3IaQhIwx8n5nSzPLJl0IRWD1OkLzAoowivCmYsioJ0hOWYgqf6jpoPQyuePeT0gaUrD
YnjXGnV8e96sNEzoN9mjcsXjEPi/KyzV6tTeb0ZyB2D5dk/h5cjV8zzlonGrRdE0zw/RL78OCrQR
r0fZ7w3dANzAHYAEBvrW8FY+z9r/lH6AiZX/tKjYW2EeQ8mUJrRBOEaWhyOOqTgHyTJqxhrG/IDm
VNcOUWCTlNJ0tKkblLNmSpHlaClW+C3UQOF8QsTibdiN/Dev0n+nnyMBAC77rqG3X8TFHpZ38k9d
Bmd/IK6EqxeLvs5S7QB7X0Nws0MKeHJbMdN4XuiJWEGWw2xWqjrm+GZlCFvys1vBWqYLJZk/Qb0J
15+MJsB4Zh+oOMY4SqbOo/dKc3yyDq+tWCysRcyZclQTgirScegV8eQUb7DPVEMzU+vjHmXqXy43
WkIz4WbIlZ8icICTqOwj5zyv0Badn5LKEeA5rfouWELsvtC1hHMLpPskfDTEzv40+s+FBV9klQE+
OOLmRfQdVRIy3OKiJTCz0+S6mQCoulsf5UYThGNqm++Wat14e7CnsnDuPvnGaM0J/x5EtCvXHIu6
HnF/wD188l8/r6unGkXlOp1MzcqioCuePBCnpArdw7KqM3349BYFs/K0wWulMAorC2yapvWSLhxc
ohggSeOKQrhvGrV+nt/4bJS20xx2djH4H1+JvXzLr14AIGoXbRR/9KG3XZCBVXauMh6EwZISt3nv
ozEm1W1on2VgxQ12RlHVIawjwxbjqu4bphfgP/fkQtqeFQaClJZwNIuWZksSsPD7wHH23OI8bFXF
NVOApR/y7vxnynoE0l6D9mLpljnJuqG+Z/G7Je0SQ7ua/oLgS3x90wJlllFIsqW+O9LOZb+MMPE/
yStM+v6lbVJjEK0E5Krvj/6tZrrJ1z+5LRJ/RpfO2u4+/J4w0lphMrJWQpBeiMwVY24lSmJsf4ab
XWyVHsSpyDrOPz8pq7LBB6lDENDcGWBgnX6SsEcsFKfYkMITL2bC7r+xJI4n89NMXInK3PFN0PmB
iLgR/JfzjLEGcElsneo14XiTUk+30al8DusGw431KBlZ14fVtOBofeUl7wok0rmnTF0Jwj1GZgTS
SUCxvGJNdjMfsqOpnoV13OySIFdq3L/Q+HWIU3CAknxQWHIYckuFCZ8AZlj+Owaiu3RWR2LXZi8C
iog3+AG5nHurEYVjqvlvcAcWB259TJDfqZxFTho8wCQ+Xi7FNVozDYj8e/l1whFw9utVa4YxRbsZ
dPpkaoEEwH1yWB0XZFucLZDGYS24vtKpp3dBuYKDGmQ3nHSgYLzGLovWhnvaRB/ZjdtWi2VzoDmE
iKerw4nPYz8SVTOs4GCOhQEOYiRAwdtmN5rMEA9nsa9RXC5kkZsHXCI5By5wivrqxdPUgiT0mi/k
yIuoHpfBKjPGk0WRTOXwHv/nefv1UyNDaj2SskTLCT9OZq3ydxAKAi99v93eHuuM21z+sZfopaFj
WFBzmY9/BoPVt76/gA/L2uzBSyalVvoAkJhp982mFiOnnnN8l2IUoK4HZLNPjEfrQ4X5Uc5C3eEQ
tKemhJ1nNGuVdISzyPDTlV6CyQnCpQmrXX98ALyBElLP2h0xSmem3IvpBXwh3Ng6POCTjm+P3s3r
4kjDeiuCOZmPT9CqIoepjsYUSlBRWrBhmaupvQ05qptxj02YnspZ+gG3vYfgc3ZaivJxJKyOhmEs
rsnfJTtRwT8F4jpTKqeCtYuJCXacY/S97cOIgTn1oUZ4cuc3o1tLvdP60d2IJcwWhNQab9SqRTJ+
AvSOWIDmJLESeiDZzLlM7PJIi5xlN1wwknx38B72LgndG48BKtn96H5B/ylk3e/DE2DV8pRMH5oH
jbn42nShFqM4Ueen/+xdH88BC6CaBKVZJ4WKzrYjYVfDNV6odnQqdcar4ftEdZDpRMe6O1JXWFGd
+EUf+GVbXYQ5hVQOOs4c5ONe7Si8ULs8R4j2LEBZaFTjYWldHqqAPMmptWzkhAlcSLmsn0ve6y8f
sBR8h2Rs0bP49i9SyWOgAaru7+A90uFUg3SfmY182BW8Y3hWIZsgdJnNBaBv65Uynett6k9ZIJ78
jl3mfnREy2ZIh4X2/+TXwPCFmnyB7iV2ba8YnDdnuf7FlEn69C1lNohsMzIMCs1J6M6w9iUp83u2
jfRLkYSP9vzK3GXRZ5/9H+SzkcQKdbIZcBSw4IBulxz0r/htvXdweqW14jr51Vy/OGUYMb8yXsJ+
glXLMEOabl8rzKm9ww9o9ElrD7BkXxkEHLCnFaRaPcPqSPhvWyqGbavv+pvKXvHZwPMKsdcYoNR4
BYdS/tr/79UVApJpSKx2thvMJIfq8tbxl5vZq4eCGHQw/gXZV1PClbbKsIycUhD4cAYN9c7vyBji
uN307YSpkYtQtFzx/lluYtzYwkgfJfyCzBKkxukQdCb3xHNA4DFl6QJjQUw7DXfc73Pt8Ij7uWW6
smt//OS+2hpZGQwNCpl0HU3jW+/0K9EqPTozn/kOX6smly8vtmTHay8zLq8CLqQtac3ipGjUk9H/
vfvL1ldqIFG5GpJ2zqxxRpvKzX45M6w+Us/w5UAg/CMW9DAZ6GxoxXcFKTqsRH85QogDbdTXhffa
U09UAdJupYPqH/vKXkOead1BWSiak1P2wUu4u+Nhj1D1CXmZLWdcw9veN+pJx2IoNCYCQ5+Pxi5Y
jC9eIJG97ZNBtqkQNHVHUG43Sdq9L+if8nAnacDEcIi2JgnKub7swRq/dddkXVup6tuWjzlY7zkw
3uA6T8Q4kbXBI/ED+yW1HsionXwOO/7Yw/U3t6SSu0ty6wg7zpg3WaYhUfwhrM4PKMcnW1Bydb3j
muSliDUjpqr2TLfZbI6Ax9KjynYjJpUnwGDo9yK41YKonUngGXqUoufQJyRchsOqZAUBbRec+bbc
OzcD/94krGS5aSW7j0zavbbCbrGqp9gpi39/dJLqwv7mAGql9OoRB+uAU0TNUb5Hxmpqj4tIkr5Y
yxLbB7ybwXxNCYS5m6HVsoNm5KZHTORHCzjH89UKb2ozPYl1t+QhOVUDhDm7BoD+6CUxldSn+Lab
1RZ2M0oORAZbeYWZt250aAss6nvIzmEl24WQ4Je0NQI25rkvIBR+EMYCQkIHVVByPF30dLfiUjgx
o8WwzOtG7EjDpMDwi0lU+/9WkSP1PyUytv6Fx0IxnS3DKSEL19cNx0Nk2if4ZPQQaDU08vFsMkor
U+4cNFDZggLgacHc+90YCRRAYueW5nHEyqiwgvVS5SrHeMaZju4W7ZTVQ3yi2IMVaCy/9b8w9r33
Ce3a5Ip0BjQMkJebuQ7hZJCEPNUgF/Ei2C8Csm5PAOJrWQPJS/YIxuiN3HODx7DjGLu2IWGGUxeT
6iOiPsmb26UX+LaaF1+DIoHslFH/ECLNZVuVvfa+zbbiUS4tCepJUxgidW+8AUXq+u9eg7H5zJN0
XovSLuwjMTet8o5vvlZ9RUD6LDmbB/6AATgUBDH5gI1avNBXgKdVTs+UV+VcZcR6VZS5Zar4Ggqb
MpVjNzO+zCMh4UPIntVjJTl8Gm1cohRfgEH3Xo+rPaAkZ23voiKtp26b4qJDaEJ2W36KD3j0/nQG
4GgQqmdXcdz4Sx1Pi78K8VymeNHZprGn/KiRRW7IYYF4NA19g9I+k+zHr1OUpOToQpdRKTApP5xz
L63Q4UzyKG6avy0x2WnwdzcuHWTrdN7rhUm5gw4h6vMuuwOY4w0sXD5uvm2RU7VlaAR/4yF/g8Yv
YCT6QFW7kdAsd8skRVghSNjorna33e1ZTMsZV2G3qqYupgj1GQ+HjaqY1UZd8++ZhWK8Hx1wk4Zi
wkf4VmwnhNm/dDOAEI4SqfdlvONllVbbx37/d2hfCQLF792ghjgcRkcSyk8FMFM0523NqkwySYtz
OL118GJb9N4by5xch3Gy9UNcg8mXni03m5rEkSU7DkOsogQgAiHJiah3FgrHSZUOn5212ag891mV
zTrVhZgvKYGVdXrAi7+DB9NzJ5ii6HmT48yQgk9fLnZddI2NZH/XwxY4AJySZK/nRGlkC57gmuNo
JZ9gN7qH6O/SqG/lllNPVWJphbu1tzMQGz8e/AH5nvGE6z1AUbVyDj2PSZk+jItTv/BIEaIlGAFs
5rgcvCAVyruA5xpCZ7Qf5Lj1pZcYR6yh1Yxtgt0Zum1DBD1UTVLMsUYkDoWn19D8EkZYHrELWCPL
tcjs5ux/Vhj8ix5dqcc3WZVpjFzi2OMrMoAFV7b6lXanR9jq/+WRzH3RL/yN/jjeMHv55MqFcY9E
czEwgRJo00Te/prEvEuDsw9NsBQMp7J6c5SD7B1Ios/2081CiWJCiDdDC2rGaWP83WCiy//zzG8j
Tec1N/oNtA+XoSSyKeCK/HmxhIdmTLir88+P6t7s73guFG7BSxhlTLuBdbKwmxSVAd0rbOzXMQ1J
SZ1J8HYqHjc1wG96V2RfY+fD2ytgMul1tNX9VT2o4/MWixoij/e2QaCSnykpHInTqIsJFEx7Pk5X
0N+tjlTukAhGWXqnOu1R9qBxuDFDM1jRyxH8Mkh7EYNC5srnlySmu2AXdkAUeC3Hwr4lITF2r30f
l3lSKSAYeYrPYLtII9WGGQvTNvXvfhy3zMnVIrHLSZl7Y7xtDenffrXn48AdjsBMAacU2hFNJ+Gu
Pe2ihn5RSw71TRKngfqGjYnE/6sUd0X1GqX0/wkSiwuhtrrz5fr2ENhPoPzoYp/08FwScAXT2VG7
3tMkA/4c/HvhZazpy5Em2axUP2n0t1kStTMiMz5wCQf87/9B1YELdhuNH15IR23+S7rFinQgmGGE
BLDSAX8Wqm1gWZkzYMJMD25Ou46FmbmYdkLIG4DwvR8QWHebCGkowOcTBl0BG7IMaPXcuJhK1/nB
wNnvKoV04XorY49kzIdgTQcKHzkP0uE1vbHigdyab5rf01DrecVoFfDZ8N4aNwRJervj1gw36yKu
9VioIpGda/Ir4aTkp0Zs6nv5gp9OwSGfMxHZnBqgc7xFyR2ngkyz2OW6Ra+dkxXEqy9uELIQN2Yn
HxfwJJuWyqhPApetK9XV/SnVInp9i2EmjOGmNxOxoKeGcgbwCndmQ4EJuSYnHxFfsFYfCPs5aYjy
jyT05bXEIAyz0dzjJpNtq+cptPmuQwKvznuMuAJ7F5U9tRWiPODr1PYia3jNdQFphCGXqhcpSp6g
oSgNyjPMTBAGAFOxq+JZbii5jvMa3CwKF+8VNEIsT30XKCOWSmC5Rtv00UJQFTDdd1qwt80NhLge
lMImzKm5hcqfXyhZn4PvWtJtTZA7lJWr+nT1KunfDbzJJag8fqsmozIJSPgNskstyCar0+Jk3+LA
vVyZh9+Ba/aKwakzRv1/t7d60azIBhp/4mGb8wy/Wsmnet94d4RRW7/CljhklaoesV704AIfHnhS
I4xAh/yipxFV6d7q+9lgL96AVBCecNoHC3/yqwGgiWFXpZmiBiJ/k2+TTmWssQ8NzjDG+gFkfFnc
l489UHCzoTDEfDOq9/u/lavxSmq5Ln97RElDwZ8ISA+131AdjhleiSIbnzElPa8s9xfXna8lvywl
b8zMkCBmjWlDT8dVcRL7JPTBkXtUSPGyZ55uwzAknaRVAbtLIkhoGuMwwiXFs3DykEYhe3J0SrXH
FeY4kVwE7xY8cgitR9rGlofnRLV4/cfGf6jF5N9WKw+pvnEiZ5aTDXkvpi6lIe/Wyv5kB2riTeOi
Ac/3zeAB2P7enxMKY4l2SNCftw/4k7zUFD4m+bpxfryUCW7a9VaF+1xf0QzExnPh8bgdHyn3h0Il
Ds5G3wXjBYMsEu6JUuE/0d05P9jmC26agPor6l/pVCgBUcpiQHm8Z/xE+5eZx2uUYiuHlNW5kag1
fWfmauZO72yI17iy45BdR++gfgl8IrG9B3OTilSSrrL0ccAVocX06uhSQ0Uf89NN9asdiR9SzFW/
E+ImPPuI7uqvXECCsPte2x4tfP1RARW6lHX1Lv9hmOJ2BlcCK+976UKa469LoFo4go6LYQ7/0eAY
3wdsXeWKjbKTG5E8dwZ/r5xMUFdSG9ECGvxNsxjvJ4HxlN5WDou8l7y4SFKtpnUVcPMtgTZcA0gL
CfVyqNPUn4pOnOAS0HVMTAp5vc4aCF78wE1bYTuL7CbHQe5sIbj6TMOBv5EbQ0hrFhXnw1xdMZ6Y
PxDhRLO86rDmZmMIqfeIHUyWtylijxSkv5qkkT2hrGeAD/7H2CEz6fKTv41YyKAfemXhwXLkRy9c
DYm00QW3EXV+0C29BOkjtAk/lkVsYwPyKx6bnb2kbX39G3lo2kvO/h4XK2br2qSmU34i+sfmiX+y
gHFhI53ek2grO3e15yzosNL0wDUDbkgQevlN4wDbEWIJyUGZb7Glzh+Hus6neXzTexOQo5xZiSLk
0bljVmdC4q6yyo63lpHRDaXkEct1SUy7tRToHYsr0lA29tcAOxDCtN4SgH4eSrjB4u6E0kYKT3id
tWqQitthhGRi9JWublWT8+GiNRpSzXNmPyD1qp+b70Wx4wzPUowB23zm5McenQBXBfzV0qnjjrrh
XoV15bFSIfMTx3rdeWHlCRXzPo9V9Beo5Oy3Iu2mFfCO5Z2VXr4ZKhwR9MHUghF1DObFUt3sC4BW
1a2YacGKjhbFx5CiQOqVMy2EAoS61gFlIj0qoQm4/Z4S7TmMhYi5Mff2GgjcInyGn/GE7e+tvqff
2/hxzxHR1akH37j7tD6W8r70VSCukwQU+WeCGz0ctY7WRxRupmN1C8aapddTJXokuy2h76qyEy0+
PoHiaSJ0+aFRpLM1rqcJlaxWfWh/DjOJpd9kP1qn5DhUXm+QOGOD+My9APHeX7jG0lfYk7Rp2KHr
z0ULblSe8ZP5g8awXUUEBth7t6x1sqQA4UVjwgX0mPbkjIZ5vqq89EEtbkf6I1odmRZP9tS8ePaV
9JJo8H4skLt19bKl9w5b989t0FtXqteLsOFmUHOUhsxywwoBr1GB+lr86oZjBIGtwzk8k8H+bfTU
IbyRvg1aNw0tdkXsEw3nOdODgRLWfRqSJLo9qTeenRAFCG9tC4RnuZyUuNOdmYxYIJ7eVuZyryoy
eKgk9dDs7flK616GTYmF4bdshnyjQGkR100DpFJtG4ixHyoA8mDtQ9fdsQShw64gwrxaonl6Bn0i
nI6CcrVVwgtfXpM4KbyFmrqMfWj780zjqW2/pSCAMs/A8BhlKN6arfEiGtwWmc/ZJzWKa7iOoJqg
6lK4ZmNJCkGL/kJGMWTgpWCqEMTvoh6SsUe7wufK+MDjPSl0rftG6RacogFWFmJbif4K1YWyJazB
WjfpJMdUifDV0E1OuHA1jgOGOxy8HOFaZrrgZuJuGwHKPeG4vtH2OQQLw+aIQsq7OLxDvCpDzGEi
ljFD/N4/JRhw0p2pCy2nJJKv4D417QL6Iin2cnHb8FfxDZKr9BtQW9xez+Z1y7Dmvltw/HQnCNnc
12Gc0koy2JwH770lOPuOR0Q4INJIBqO7Y1tSxhqFEsamXEjWjOXaCGLlBVTQ3eBrlRKtycYes3Nk
ey1eDY2Wk82G5qS496+nurt9t3zwAk3opvLel0J72jglqZetCWZRMXKDhfgH93ayt5CtNzyhCJLd
ASpMFIxCt+GL/7fXu6O4grfss4q69PrC6GuNq5Y+WlsVVQz3VYFgaiLbpGtOoX1t7qMor03JQ37N
H0Uh3tz4pKf6rsR7kusUvynn0nuJY+P/SxnXUQ3pLga8qQYJlJr8PAalEUdYHjidyu1zzEVAopBC
qp+hQzYKZ8YPsRcJYBp4xNZVlND9SBgzRGewqpcACPeqKXg9PUQohXjt7C5FzQBIqcLu9B/mzX1M
k2lWqnMvZ5sJiGrfozi1HaCLnbZPk4l5TbhBQ3jFTjRe9s7KwbuuW7T28O9+3ab+RGHsQg/umLqy
VyWWjmfCxMmQgi3n+/+kmyrAI/CB2i/p+WrsrJi7rx/ELHGbdUN9gwKwHu9RcRrtZzE5eGToFgky
0SMdIjbAGSHyb8XKBznLEOfVae5A2m7PgmLKkU68EqfeH4hfehnDea56XuYbRvbpWTY6WukGojgT
R9M9EEko0HYuHXqwFfdT9aNTkM0YGDCBZtnC/nJVhacVbJpxzEgt0HX9IDAHvs0nulYsVQe3xjYd
FkzXukOybAKHKuZ2AHvrQ0zqcqWgG0IVis97Ml3y2makpaN3zdoMTXTIBDOWvoHK24KDZfq4iCb1
HnH8oj/L1zNArfNHBlfu6YrUdythq0dFhq1dcSoZMSxAAWgRZ3vAUe38H2yNrPNPXEiu/9AtjwJt
JBivFz+DkTZLzyfIJfjFo/s+69v80KHnSYkQwjOeRquQG4ubYTnsxup3aUX0Pu+clyz0JCmsprdj
JpcixPWfcjXYNMLnZ6aY4EuXYuX3e9B7fI47PxqTuKfqtouLUHaaO7t6ggT1eHJ2e9CpTyFvKdTX
w1o9kisIv6obOR6kBXk2a1vPiVgKHHvLQhmsttc1HxV9dAQdfm4CJRt7EBMiXDnw1QAcnj/H/wz8
7Jm0xGofu2SoXjmNbqtcE8nX8aYRXSgJ0eJ0hA7Ed0n3fRPR5/RYtAhVIpsHNMh4qEwZlQ3zWLGE
vVphkK2+8QG8iKkYMd1BhfRrAR0ZCpcmxHc1IiUMV1Luqwx81d9Tt+yx5T2pi+I+iQTknkA2x2q2
am5/kCYBp6ECy5MpjWTT+1twFWATai72OU3awQTogdXg3BBGtMrbYI5tGkfxKE2kjV8u1FnSWgCf
F+Sad6PK7YXEN0hlVswOgmVjOB8lQfkEg6gagFxE3zIJbQjI6iDodEE4rzRg42z840P6A6AR3ZHy
gTxU+nr8L8z6cURemPWeNHE4wqpIMYactojrFtETOkPkIXrsqt6lAS0QMYM4gB9m2wGvHvh7dUmn
Mv2KnpxUekK+jANHXb5aA+jZqzrnCngXgXB9E1bzjQwbt/7y+0vOc2x7Qqp6FCYHmq3Ved+LMmvX
WIaaTtVGLE/PzsSRdZN1bNm6d4/8pzYpKBzR27hATDvn/y61wLEH08OTRQStXSS6huwhYAN6HUtI
StmVcHczGUfNddDF0IkVf170UJ9zrHSGxWypOZu+2aoHRtfB/XcFLXeTzSwA9Hh5mYhSYMqardDG
UaGkUk08+dgq92x5iLJhFMpdAKwVzHJCAWLjeAH9H2rleGWHhRPkAjGsjzbYFPdWQLSK4TuBzIIp
MpnvOIe+KLX4n9IOjIBGqeoCXVAthbjPEfNJ+evHH2PemWSaf0LuNjUWl6s3uxNWaN8iTj6SRwi/
bwrBuotXYdaV/w/bRzxfgapEq/MXjOM2kUcwU8Ajd2gm2EcvkS2G0Z0PktHoi0/fTURwFXQvuit3
ftByWqdiaTiphmoe228C3UhjCp0KUtZsj00PurPrR6CnA2hk8BxLIcB4BHYZM0sepPn5jpq72kzC
ka5K4I4T29E7MOd85N+QFuN/gqUbNDJwk8ftrbxaP5mU61uNbz7aAdilpUafwF3dyLGuyKupHZTS
71Q9a2sviFsI7UgMQEyre0YYulAjLbuCn7h1l/XGXQIXnfksYL3elg9gPTNiWhfG5rZU5bPZUkG/
M7jtm9WJEwABLPut9OBKIqncBtSDqrxYizkkbHQd5a9vNg4nXRPsRNlTqj1oL2LiKEKIDpzlGjPa
4wdV+0a3CuLamkQ/FDfdfbreVhx6stYRcLhLI/JD4VD5SFbhwVZVGHrWgaxZUgYLfjABY1KHMoaH
VrJnjGoBaydkgHYz9FxShYjRhOnY55oFXYWfVKU7aMgRS+E9KPIfD96oMxEwKx6pEnsC2IwT2Kfz
v/+wMT5cgSEY/oDxQZaLRihNcJ6pRR+BZor4vUkKdqyV++napfQ70cHM+aHkNQFjRcQkkNSp12ki
FEq9K6308MP4pkgqiO2qR6+/121DiChCP38BygMUqwILFeqTYcd3Ji/9T1pzQwAUbarCzjAhl1AF
CPs/eUvktePWdSi8YYSU5RCaG7PdiU0o/5bI1BPC58zGRVs8unX9WKygPhEIfjuF/RGZY28J9Iiu
MVFAY0kEh1gw88gMdU3kvCBZyOoKG02ShXv/FXHAv9H1EFbSx+cISHvoqxuAbxMezv7mpp22l5SR
bEmUNdY/MY3S6o8PjDEWm7JJqe8hWF9QkS5kOQ12pMgXFfaJLqiVGiNld/Z8+r24OXh8uBBdcPx+
Xmvdf88ud9R8zbc/osCdXSCX4b7bh4FTL80I1HlfjDNV2DmQ/wxtF+/aVhYkgmq2QuUMzmEKlwn+
r+dCVcXOC6Q1A7Ia77sQibDXwFt74VQOD2O8G9wVQczoBnn925h9oBUZaKyed0QZ0FiWBHMjcljH
l4afN3NSeFnNeBUytSTGeOVXsoHLSGP79/8EXxl0EmgYsbQQKf38mapg+XT1niAfKWAUzPXRNqt+
VZNuy21l8vlKCHEEJ7WUj95XbSKxwg9j3NxunUnBYZX+Zpk8Xb2XcWOlDJd6BfcEkIxrmspi860D
E3cR2m+TNwt2Sq3OPjLAct4wntk705gmX3gPjm4HFQJsA9KpcViiI+9RZeUewuNRnl+FPPeOZVf5
GgUIYTGw7ZHWdeITZOTMwmSeCNqi6xaozhqpNGmxB8+QLt2kCE/W4yofacRs7ukcjypEYmnW99fp
1j0pxrmgXQaSFkIx4v+4loS+znI+6iPru546kK3us8oB9qdwx9Ifl1qAF1DUZzB3J0hOmaxgLFGJ
PgAZ01i34nGRmNK1IJnAwzRqUBpBqwnceUGAMyWLkRj6qDY5niKhZobLz5fQvBwRUN//Xb2vsJ21
ev7s1X+AM0lv7BWhKmrkMeY4hJQIjviiNE/GJWx3baMEKQ4bBwmSDPRyOyATmSyV6Pkxx/YNjckh
1h0TnKptK8hmnpGwQZvxYH3sSsb4xrGX7zYmQu9o9sDI6EAM0NrO0n3007Wl0mhlerCStoOFKauM
H+NEN0Lk5sWGgHIGM/FYY2aZHk1wOVHECd/uGIqAgIUF1gFwld8nTBcWOvmljJ183YjHxqLJST3b
LgQZ9B3zlmkrUd0Xy/VKo2KNcpjqT96HNQQqV7jYxM3ARnbgnLwc84uM+WoeZ68wl0rNhKgkagZR
da4vtCFjoj/3PBLSVnN60MHvH6gJReMI5PrWZR55z1DI2zy2lYEXX6CHsWBmjiwt4W+qzsxiEBCs
dVlC42kSCWAfGvz26qOwsPiDc0CuulpYqKNK8LvxFq0ATD2fVHwL7RH2hwZsaZV5hPIAupCa4xXO
VfoZ4KC07DMZnrijGuwdFixRxBCt7eVhjMovDCsjANVPT3VkiX4bnkchnnMWosIjDQt53TvWOMF3
/cN5xBPw9bb57AwGK3a47psWD+XtA76U7z+Bjv4PV8ldVDqro4VgMWVcLx7ZG+A8XB4/3Q2kY5sc
RItmYjZJGrMEMsSVz2dN74doYVDVDkcDROn4wl1s6UWAr2PLC6M7QdFjxF52KsufYquSnfW4dJxo
yMLztGuDzgylYxIbQZ3wUdIJykVlmkbjsh4GjFWQRbAgL/qP45fxVsi8KG0fF4DC1AP9qGlBOKec
GOgB4NV5pRzRgqjy9ivoAmyP0i6zSFrFHrkFdGEh3XYkL0sojCyuQ5Gqgv7oBEX3L7wVl8IUMoEG
cHxGSFg3P260yKAH8DM+Z0lUvP9E765f2LFogcgMQseEQ5OAVR4xzDoS/pc7I08/AvESdBlqTMWE
vAbIhsJl8Qhl9OHzKVG+cSQl8iCbstadNhYULdul/KCmEjIFekJp/djxSUKJ6vCRURAlun51tQDj
mU1DrfVJ05ue2V7XrB//pWL/FBD2aqlHk0fExFitIg1GjwqwW8QotBBXiainJQOsVbrVQ2C9qVBa
5tDxCdRTlQ1jZ7Xnoriz0sy9Qo3szUknTCCxEU8cIl5LJrwbhI3vPaxIBI//geJ7PtsCNceaJ4eb
dIpboh7jY24rHKqNS4mWlAAziAS20kZ2YM6wd1qrkGIul4tm23GjYGu8Zv1h1bW1gSaR3tZmC226
rK7XPP31+ToOoOa9QeRixiXZqUba5NvCql9gVCmcvukyXCrgkG5fmYGbMLaT/WuUjduPWJg2wIa+
gvRZWaRZxicz//MtSUJQMJCe7CzSM+ibR8IPjyhRlnMU9DJ9M8UDILkcMETgEpCf5q4zFeU4CKfT
NwnN1hygglPZAyPFl4NwAHuY+Rh2+DDhz0gQVrQ4dyviJxp3TquDOKo6fXqtkZpgrRAc5gH4KNg+
dfPNIPTcKfoKNeWdLse9FF0/9uhG1rEceaoM6rxPkZl99x9jSZLYaZGKv7EkeHJ9B4y3uDgmVFMd
sLKkfcWul0BFv3V93EpKuwvG+nJmk+rvZ/0+0FFpf6i/Kb5gSBxGomHwNRn5rNDx37co5FrgWz7Y
1ns1LNx2IBbBaItjXXYdgkW0/ZvcjheRaHZ4gdfTYUu5cHrKtwD3c4JA93alWla2CbcOCKXG11XW
7QIZwMZKty4lomLoONENF2YwBcBd6imGLYmcVmC+R5rGdoY8eMRsE92hiBHdfLXoRhkduPC6lYVo
91dEReH8IXGoVptmSBJuUUZ72pybMRztdogOKj6vmomHqS7GEFFHLOHhz3KgNi7GXPge13tWC8uS
iw5WXNW8ED1YB70GGrF917oXcwtIglqMY+Dk/wPcz/Z/xN0FE9iOfQWOKQzaADNY38Tu89wvYpYv
VfidPLQ4TnAF1/+dGwHG2Txm/2/0yxjdhkOIk/stSTzmIAMHmmTo3dHIO9UnYBg3oQczrGT2Lojt
ttSZyDE44VbH+zM5+zW9BuNkrd7awqIrFRXQ7xu+wZ9gef1hBlxQSTumAqQ65pL35IbpoNlgvgK/
MVNJ2ITp3Y7KhIUOVtplP6/Tla7ZcDnR0r0y6doLfhc+cQEOBumNskrj8k2etw/uIC3fVi6d/6dO
aOwx+xOmml6zsZtgxkJfARuplePWmdyCbosKFcELjA41NoVaC8X/4WqIVprWIGn7nwlXxygjb5yf
qtWBu5w4ydDxfdMOftrqlftbT56EGvqfxgBheJZMIwwXY3wh6XCD3e3sM08xS/T4l2omqOGP0vel
IqzSkbmzdaTKLyJa1mDN70S9K1ry7acHXbGnJyfOpuHutIm3efFHb6dkGsgTJIosJi26dEphlkIs
QsjfpgtxMUouIQ7IIbB38qhYx4Rnac3J3O2sMdlEqFAZE80KsdvmCZdNY0zS0Bp5bNtroV/GO6Ja
Kn6KpxTXatnU9hn8v9Pb6xO37vUp6d4hu86snY8IQSp1E3R8nokmuZJPk1QBC6Ggd+KChUz3rr8l
ydYo1J5xF7I89lpq9ZDrt+k+NPrmOkw+aI0QueM0jUcTAkgjKTo2Th36E3ipisZxfKz4IJlB5J9f
QR70WuMhlt24z3FJp1sIwr66gtZCw+HOy2BtOuhPoHtNHVxBtv+VGT944HN9mchdbLtdgezxF/XR
5R96exN2224LB9fZtMgXFIUQuxBrApZxSY5auCGyfQ35GY7kQhiRget6Pt+gl/fm4MsZ4T9U8BJd
Ykgg6zvkc4p9OS+SLLlak9sj84nzDuMi2fiZNhnYUM+xQLf401gMIN2kXpdRlwb2B8Saalf4Tmdb
Q89AWPxxInPirOd78eRC1qSk8rxmWRUD55Ba3cVjjoIqWPrdmUwc9ocG2s2EL8XF5IWs8oD+Z/WY
m7yq4eLh1Myovm2ZJ1L3ZsH28aGvOMumNOXCrirXF+cF2CUI3rNL5Ox5shTisQUteOW1Xo2OB2NA
ZYyLjBkRBd7SclRQkCelvqSRNo+hfT874cQ0YTsXIn7DaKaEeGTSYoqEBml9bJ3IIpOF0QdnBXmt
ifH91h5p78Sw4JHHIG0WNq2/oz1COMsMclkb6JQmESGfG8eOX6T/CAJWIwMUoRbxmQHOTIa5Lrxs
FwoA+lKkuPr1ga9lMKTvJ0vVxiuwH9xCO7/SD1/tSlcPOuQAsbbP/qiG+thGkSGwIc2QxsSNrIi7
ObFBITtcnz7d4ctlMR9HiON96uerstMlOckLt8AyLrfLMfEjtDGDuqB2xTbvE7mcGfTo0ZJL4iKR
1MrnBAb9upioBrmsjTfmKmTkfYszqINzrvUzAgEnJNsY9R4eEg3HM3zManU1NEb8m+fgBbsn04Hv
cANQAK7+HlvBJ+KkqX79UJHkvAcioRiMhZ1JukCyCsLRjKU7uMdivwY5j9HITi3DKQ4zbpLclMmB
DXNZM6tw4yYL6yTR8wgP0DFMmLDrlKr05+9HaAkv/i5a/GzDrVmH9a9RXn6njGS8lRP0e0eBh9hb
0w+TIRZm/igLOGbDWjK9HQbEsRSVcup2KM7g39M60P7qeaI0aOfy5yIyOOar7mUjeESAF2glqQri
E9uNCWBmW0zTMHhZFmN5tpB83RWbYkyWmBjHcHGhzFe4Sw4WEZLxWeEEdENUy6AFsXyiH6ws7jKP
v8APZ1DynEgccbUS8z2E55yW3hqYmlJhbK5gmUARseVjETVw2Nt0K3QjkTHyaq1axfSRq6xbmcI9
FkBESPpTads//8CXTfrp7fGYuCgfPAF6jWt277gfYuVPUUPsCa3ZGpGVp+NRhxrB0O1mHtTsJRmQ
w/08l6irIm7qin2fINTvCivj7e4yYKR5YkJi7zcYCfif5A5EGnEvY1Qm5Mq1k3cJp6vsz9g4klBB
vQTI/agTMFfCHwiFQHMxYjjvKh+HA4pw2ALMDXbUxWamQCYpDkP5PhNo2PMhthcZAZTSGT5BoAI4
YKIpBxdn0bH32zuimkbG7OdH9DQzGWW9u3If3MLqBIGYt4gXQlwlKsPTCOdfs25MUDDV00y1ccjr
MAirjlLjpuHRGWb1JblbF4hG+/KNrLEJX3EbhAXDikDQ/kMXV0FzryURYe5tn3qrVBkUcTtmtQq5
ACCvApafM+eKuK/Wroexjv7/oBfaYXM9RXHWjvFdci+iZw3RAF6SviP2ABSsCyb3PlJ6CJJ1AurF
NEsAKFvpvN641mdd1XBWuF71Qfhr9IQ7CvDmIBQ/4FAB/kwTZ5HI7FRGpI87b4xVK/th2GYj9w7Z
j0NopijIJ6hvyFdkPdD3EY78jj8y8X4EOEan2f2CriCs+5mxhQ1jwy/Ijs7MKHf1qC56y/7WB73b
qpLCrNiG11NZZa0FKzxrc3VSYUey8Pvb5ddtgcFHIqrYkOnvKSqumMDQMHbEdyitg51qUnhg3huU
zeBjFQxD0KXawp07TGvbg1kg89CTJ8/rGYTzdQN4Bjwug3YlJYYXfCrdaVo5f67KurCkIDYEtHiS
2GsSbOkyUQDncBc/3138wDT4xWhLfQsW+QnzOuZBGOU4N0M/MrbJfRTUP0j4Lz1VnGv0qgQ5zzNY
/9JHzpOekmxiLEUn2m+4nDxN+4H7EjwDocZFvMG+D/1FZcjk3kDXCmrqpWvNmB/BN31uExmbZHuT
fZJSi/1xNA6d0Hh1gh4DRXCtdaS2WPMRyUJi5z0vT+mu4HvJ9Eok5lTO1+kEoA3fcdXp/TQ7QxX6
zZOdtd5wdQQeuHAauzlo23bGXk3MrwYR8FhNIWXqDcr2rk/Avx6r6Aqd4HBf6qjrmv6o4V9Yz0S+
2FKxsMHpou5yvDJB9B3hLKTtl9HByAPpGKgnIpPYVg+xQx8e4+26rwVd7pcykIXofYhANIwNFrgB
Y0BucPFTJbt8NEyF7SIqeTBjvf9GGr/you2bChOXF1HE9eao8NMWcM8Sy/zPUMAIWoy4NseaDO2z
9sZualnI5aq15qPTX1n59tfXjZrtCedZNrJD7vz8DC/oeIaQwUFDYTvrpEYKMNwEv3ggnbT5nLXb
Do5YvInOXFbbB2YOGycnDCRRHX/VV0Rk3+sw2CbbOEUPutzeuwV3ciSMj4M0isdmih9WlTW4QgXQ
OjpJa2AlK2A4FmwpNNOD0iB+Gk3al3Yki1eHf6bQfIB/TQ5u+31tp2MulCFYY4fTz+c8vfbLcsdH
y3MtsnA/WnNf2Ip8Oj0kQGX7aDR6/EpqANLUiarmIRcwWnVOf1LQuje3wpVwa9ezz4OXiHujb0U8
5oEXumq8oXRGyWyZHB4vk+qB/9zboRIwsFBM04S1MnS2k+L+lb6VL10GtrT9L6EdGHVdx9DKkzU6
+4Wc1xjHwajHiqfxSw3Qn0apCP1/iEwe+YJ6XSSZYc50ajKYuYpAR7UvVV8QAnvJ9KlqPfydy5uM
jckC/7jIAfL4kcU5OdZa2tGJuTFvyRv3nWNB0pgA/lhj95OCsEt4esI2+n5aT11n8yrlhdcgLDk4
Z8649Xpz0k3nl+mcsqqWsvpigBLi9hMCyfegSGFkwUKV5gt1UBAzy/WSubohAzFhnQP1UzX+71GP
5t2Q065tvB4R6RxsPRQTqs69qcR6jqDrBPqAVVxMpI6OPlMvNSeF8BltQsf9M1o899r8Ib8PT0RY
dXlUb5tqwBf4esdxv+wNY41gGx+VfmMV9Efh1SWjLYwiiqB16tEEjwJdixIR5UPebTgac3pkzv4O
AjSZux8yD0LdJ8TagGsjS5mu0OK2L4p2pD1d4y0B0bReB5v109YPxitvjh8bGl3mCmCTh201hfzv
0HL3ql/TrVmT//UPFu6I7jBm9uX6el6mKHtszETJCKeiNp4TVZNrYGsEnzuBJE7q0XTNlHnWnjko
kAMmdnTseR9HMZndtxJWaN4bbCSbJALzvXT6lX0COcKhVV/YR+AIp9tmRjemvlJUTydpdqf3p4AN
CjgHLm0GJdDSbkSToHVGqHlD06i2iYaHD2Lput+zt/ukS6UAF2pqRdLjs0qByNEHOc6HtDT6Dw2C
mrUbAlePoByfn/bj9zy3dtkiR0TnwI21AtAj7nIRAcZAheJBxz5YTuaKavQjNJN9/Lu4sw9oxKOV
BLkDbuVXFHdzQMMx5zqbgqqiRu+b50uQQukrVGjauiCNKWTQ450y/2BNI0XMqAHdXk+QvU9Hl+qD
Bd8n687yU28bfA6lQs2V5Q24y7ibKsKX+epWXg56Za2jiIaPVS3aMDtMXmyhkfh2Ua/w0xwS/wsS
unVi80iSANICmNXDESn7slUyJ2jp374wXEeivR5+FkkwOkbxZ7iiCshwq90yPgpF6UmpBLRvuTwY
q9z6gfckporKjNLRsiBVczBBcQJV6gZpD1fDuDtzW7+0zK0/em+r+/gGhhCH7BoiiKg+BIogU9NP
z+sE3uCdcmHmjXqfjIOooh6XzQbzjTAxiRekC+O5Bg8uOrz6DNctj9PrRVipEWWYkJ/3PRvGMMlx
plreKU5STsSj98j9fUPeYws4taGayM6awNWOZl8En/T3M26QnM1dXbxVdRh3FwpYP3kHAZqPGOHz
lDBR0tn8dvqqesNkCgjEuiTQo8RB5FTzft8b3tZAMNSJT5CNsg2wGWp+9+DwrGqqVkZ6VHbdpDKc
gon4UiWHZ43giKcyxjhtRD9cw/8iRMSiJgOZuPy9oQ+keKhgGsaacJFOowP6kgd8OTYPPPkNyOpM
fEXj9UbzJ8o/06IEdD8DyalaL+zE10SRoPOBvyl5KwTOzuJwB4dxAWattreRCzAY6cuM5r4U0Oxg
XJI8OxwzbfPkr8bM9F5/abU7OKdBnkopttw2RjfbfC2i9lCrtpXKweZ3AhI2SbtMxtC/Z6Rx2Rbv
NSNOdqvc9zCNHYc1FrhLXyyzM4j4Nkj0f9Hl5jk9TKSGYHxQTOaifcP+xy6tO8JWFRfjWpXpDvhO
ICfN3IUPzZ9jTxir+Gy7T/UTMErG6KBnFlh5JpR84vd3nnXiR2zB5Gf69/HQPOHT4E/FBSidCJnW
CxifZEUXWBJlAX3T3mflDr8/QWfKFvf0ks3ivbopO21oGMyc3miAq8t7oLfBBbpMIcfdqtchZPHk
2caqvE7qSu7prF+RGV89r9OXTem1quOR+ASM78z5OLeCYMTFAR0KdWbs5LDDQhmOxOj5blmlARMl
R5Y8BgU4PcxFYWgCRdCPA8AOGv9KaAY0EJBWzBiFctMfqGbeHznDuO+T+tYi//Tcw2npLf1k34zu
nbW8woZVQuyVYkh9WuAM2mrOQvWiL0aKe6ntCwUJXbMWofE/FrvKRPUUm9Fuv5EezY7rmfL7UsZX
lensW1n3vFsUrHMYybIzIUqXhSUUw/5LpDdKJlo3zDJjGUdOzu9svUNH0aL0ly3Db4PvxElQhzcy
kh+Lp59fJp00lWgvu7AGjniTkxQwNMi1uydDllcTOsCB+rUGPyYmzxSpRz9uq43P7tSf4yxXAySC
yGwVK4urgUJ5/e6rE4F6euGU35ULnrITgjqDfnVRr7L+Kd8ZiTwg4j/SAKt64i7NUOsgQdSP8eM4
ZPEtqWOmanv/RGFRxlVmCH8HbBoW2blCgf+Evwe3VcoGSohITLZ6LzBL5iN8HX3ra0+mpE0CVzN9
lbmEBNUVxvK5HFq3BRKHjRoNimoezb2Q/iS4ERB2ooLUP2C9nhF4Xp84bTPXMctyI9qoIB8n/vMA
L3uPG1JKZzeTZzKPb5F5fi9pG8/3yAXxd2ATkb9YLP7DrnNcHxwxAEJlRFBI9pD/twUQpgV/APDs
VVKcuIq54QG+BlP9EcU8i2DuCFFbe6sAluiRUAjrbRAGNehQvlZNjp15KhWSSqLnDKcyYV4qhksa
1ySuXcnUnDduhsKYCp2KaQJ+uLpLPlm1hF58KbXPrwS8gBO6imTcqXBCw3TLfjcYw91VZThBQBA/
B8G0KZw/OB2PU7h5VrCMaNuUSC6fiF1dGoHOpNwKkiPZNXKFIPtiLqoW+DBu9gjSvD7biZUwoHp/
LwKdiyxL+d91n1oMrqOQwMWkkRe//bdQRKuL3Ks30u+rtnXWX2+1bH1De+EYtlITa5YvluT9AJfj
KZAHL3yR0krZf3kejcnPR6SOB9HmIhcBnX3GjYlsyVaGRFBS7cIxHOIb80kXSF4m3QfmFS16ZLlI
gXV9BgsJfMPTRGC4/YsUTg97uzo98ioSJS/l5kySbLuduTdK7hHwA/JP4ltA0U8qtOAtgKEL2m6b
wmgW+tIwWyLcDTS4TJ/DGXWfHfEUKCbORAGpDaQFlWAOI4vy+4Ai5kMjKBtjun2RkY5dHZC09u/X
Nq1AWFmEjgj1S4Kml5si8ROOmYBvup0fcE1lxBUmLSNmWSCuCI6Gvfc5dTYJ8OLNF74oSYAJzKov
5nCE7+yhb/hr3c7+xvPjWLTjKkMcPITvgOBCqhTyDrEkZScy4j8Dkz46m5DQQ0lbQ0N6A8rjmOOI
0Mku+s4fYliD0OQ3L0nrdrseic1+wtTUOJzhAZuPS+v1sLZY0au62zhmBRjuAnqLko3hsp52oFPD
EEEafk5LIpGrAu76qK99RJ8nS3ShIvNCj0cP8F/dFUvq4tHDjNdFDVHW+sy/wZqw0n3e/Wnvl8tw
f3WPWgc2QtEjbvDIKvOC34olkGS2wNVmJhbqdNzsp/An3wYNYZbEKIMLxl55qhRqXzXsDAT3IxnT
VSs3Dp18Ii+QshUwBZB1qGZx7Y0epCjZEQxH3XWrol9gLvIy8knvKFDHrO4haXqqJMxKjjEgOnMI
f+A1hRJdlvV+q7ogUJnfQeYPXXn0Kx/aQUjXEAfHozzqoYB+9ib8NfM2Rh+wLIoNKKJb65U1iMM9
/VnodDvrnPRZTfgVlDIz/s7k1xJGePDt1ngaMsJPh6anHiaBA0QxWNQSLTYFK3IkTajxBS9c7kxb
pC2zCCOqEJ1d8bVthfQJ43gNLdHKDQBwZrhEV0g/BAgGva8Le6rsmYgdXMmY2cV/ELDd/Z9agr6j
gbH4R5LYLFSIQIjV0ipGv/FGksidLpYR+tXKK+9s5FFOmhF17XsR/UFkz7e/oM+7exUHLkON4Yk2
a3/uzduQtuBJGZZt4wG3awW1xKUST5XoHJozIetq44lrgw5B+iv2k6Cenhhqtn2nNX4DOsEfiRXl
hMpUBBbJZr8WifuCdKM7v4LARRdWRqYYrKANwb2j5OtNuDcUeRCqA0uqSTdCcVd2Z4TN3KhizDDm
vD0XbLnH/gnSBYNjQPEeJx79JgBTWlR7JumKjiyr83DtTW53gQsfEnPNmiBU+IVQhCIvTFSipbgW
D5XsSrGrJAoO6/vnxQG8lLDkBWbmZdlOTboSxg++TXrsVkb4jzRDKRXH7R5at2nnGchSxKAiUCpO
e2PopvwrRY4mirpIeqULOrKC3JEIHzXZDQebbynOCOrrCoYO69skl7ys3aU46mAyTChLHsaGL7JP
V7sL5cBWMy9WVgXYn4oXDMMlLQpv1Dmxan4DAYlrLSFuDR2bSiG1lvemywpT0R4huOGr2WoLYjxQ
pfwgkHyKiyRPWEnPCIFyZA8wWAY53W8FaYbu0U0FMd8SMSIvwNcGp8MP6NCLnlhL4qvyHe46F6Vt
mCml8xNSIERJVWk5j4eGAAnKDGm4O/PReVyPNfpg2aPbqtvN5tv4xQ4kzZLi0n2Eu8Xwwnxos2/d
5/Q9q2ZWll+QLfvljUa6xpOpEujrugAMFMlWkEiWzQhGkB+BK70Y2ZS+QGZGiRNyVidKyTYxSVW8
ncAT2No1qXtqQusmp9GnX1E6TC5w6cGZBlAn7ir+9DwHq4Fwnp9ptS1rL1pC43VHZWH4jtzjuQ+2
f2xGWjkm9IvSN2N1NmQ8mNnfxxoAMWZ2TLsWGhP9XoGrCgmfYeoLjbrsGE7J5aUQQXtZ8fUQSd6H
XU//DgtNTvQMPglkl1STGsYbNBvnvTNXa1vcGhy1d52Aw+7Toh/rCeaTVFLfzPqgHvi3EFOYKNZN
7WiXo34cGOqTTkaImXKFIl6JdVD/Sj52LhBjb3SJFtNPw1mrDgkykqZNpQzIizfvQ49pcG3F21dE
QZAJ7ObsfwcD1DBRVXZi5HHcmaQB3nRAllrrLT4pbl+NRZVuVobEkzmJ3xqMFyUJGyLTdYrdk5pb
USf80GZ2lde40+Yq3p396Dww08fYhU519RqilZLGmpMXCvG0pT4nsCuTQQm54E0ju/fDj80mjT3z
nyu/lm54uAITRsZEsQ1mmJhBcT0V/wSEAoqPKAVtroZl8+GWf+jlJwrW01b+2/Q/iSMiDRX3dVaU
zTwlpHCMRhMFLHQWSOfIP8CKWRPuJ3qs0vZmgtTHrNhN7BcTMRxoBTrSO3+Zf7+/YgTdaF9MfSY3
dslCg0YW5Hatkqv4Og6nvuNpA7c9wz4eLKE2OT7ecAmG8aOFXLBvtMspVRRCbmX9eau0Ip5RjpIF
7SrU3fONJk0ZTO8F7YopXmjiy6GxMkyaSbia+gGbhoFYNu6exCKE9Eoz5ZdNAD6MDNZ4tdbOjzVC
Wq4tCRTsGOKR/GvRFxHgiGEliZlqmucfIdSRyYdij/QdHvDXcbphdCqatHAMtEKwT1NvYhfCRLcN
MLZHhlfDOMm+BwivMelCG1uN9XdNpAzsDzH8uHwxqhkuoR8vqklTZEXxi+y2NF/I+bIbv7LXr+u7
V4BDsUW5/5qYupCXlG+Xq3rc1XI7GekRmqm+Un/MRzG2Lu9Bte77050uP0zfAMq25QsjeDEkKMm0
EPm+EAEEhyptNRcRXfUIlTgKLFUmm1wY/cZ+5+/3OFqAAWu4C74dKq80D3i39ctQBe85dHebmUTQ
8WU48TXNblG7hwlTv1zxHffBHVGZbOJhMM1WeeQpviDNW3Lg2gXsjdD4A0Q25Yu/1wTMjtX2aegC
CLIeqJQF6kDI5iRLDGf+VGf25s4K9r4GWMN71CvVTbHWFS4CZDu/IIVaDZfRrz5Xh4BHpOnAvLoN
aY4OdH7RUidd/GNW3cBWrRVDgo6eGd8sngQDkkpv3sx0jOjvv9oi6+luLU2HzSuxqS9uNrxGfSkR
Qwea1BIVwLk/XsDDpCrsoyOhm5LYiWZZV/5Sa+BZkvA1MbsmDgacNc3ajIWKEMshN0ecE3O4V6Ei
+lsDNE/A848GXt0Wkz3k7zNOhWrBBts3Po0smTexpDTQIfqPPhjcjeUBlkgA0/9+wIPlC99USMpi
NuY2YNQpvkQqLwXKu3uFOjqtZS8w2HjJGcw5+iKpNBE+RYvxYk7s/vFExzRHIW3N85n3uoR3xrkj
gzQpaCbajIbiFhR4IW7F8ry21kjBHR8QqH8w5xCNMCSe0bZjQhcjzT2LEgSVdCZDme1FLIv6Lkn6
jlWqJ/b/mhLMg28I4KAzvFDRPAHfRBmJ65sZS8ByGbiRaCjuTA1VeTGnlKLrWnxP/y6iTscZFA0v
9sB8IED5KN12qoZHWy27syEX9fTpCmc5T1SYvO1aQLDVzgCNqJVLWN3pwfI9NWRNgavrIO6Nko1o
/m4gm/JDudEpT6A8+qCAja7vUaB3ne3krBLx/PMUjLvLfLCfMEMFlDtcVbEv5WaY9AH+kcsVhjSb
YMarD6eISHtwUSJDRYcmeYBHk5wWojZ8yZDx0RqO+6p0uIZKkWdgfAhKd/nF1MFmy53H+63vIj/h
OnL7dBC1tZGfiNfIF704+KBvYrqzlty4luJ8ZB47E2I6Fe/6FFT0wGMMQqQgW4wLeRvFkeS32cBs
ZNhdwhpEHmF3ff/aqNC9H3vxTWP9GPCV3xSOjPVQg1lhIpsG3as4afk2KA+xq/p18WkR+LOmfuuX
91x8wicioBBJQdMOnPp8YL5ri2sRVR7aiTTUcLGcecxqRYZCgvEM6u8iDQjliCez/sTTjnOZmSKd
b70IVILz87sTAtWCtn92hYrR3KZGLBjg+ziYuysT5DOz9Cq2YawQCQ0OuVh5xG+hfmc6K921dZkW
am312ijG2o/U+9Mxnh0EOrVrNCvAtf3rLCyupV6Nmf8GtaQ0BDuLXqflYoltXmocY/UJ9KmIbJEu
I2vcbpuUv+PiFtDLox4VuSE+0USkH/qV6nLh6gw7uIUsdOgNxsUNXqwWVO9OSOB7CzSODFL6M0R2
RhQc2Btb98DoMxm858/soSZQMn82hdejT5PtGfekFcVyDPqVy5gTxCtoJEaSYdbAZsRGsuuQK+XM
11HrBNGOEHlD0bCwCCIKXeo/2v6Psz+Lupf2aj5J3wOCL0mc/2PGbnplwwT5GsMDDfhjNZTgsmdy
5AuDC8P++Es+iF6WdIsKQY3MJw+da4y+ShZ4sfrROwgwZimBRzfJ0edqCqWu5TUfrHKVwOoT9EU+
wWJemafG8ZEoXobbOiWeJ5AP5u5tgPza5osAX3Ub3BVRaBBpQ0aJ3dDpOu/yTPK7wd16e/xQRIQ5
CvUS7AZ/GL0n7jhZRqutIAsAaNCHJbmqwH5laPbUM9+7hT/cSwDFEtm71qxOJh+TydurpyTUcwwZ
PijfKk99qmdkn2r9vZA7lS6FPDXRT4HmwtiHZnx4YRA4ntFs/qwDzctl6vBGMRe2GwzUNClpNBvn
WHHX0bkJE5CRT3aTYoueEumltVOdY8G0ph0y1ApQ3ZlrfEGmSVrL7ccj++a6/+sya+lYLgV0Nkho
YUEbk8nhtUbhBW2muvPgjP5sfnzn9FukVcDwsXpWHYWaep3Kxey4kvsM8+IxHbOkwRdZmLIGRYpC
zq2Gp5xqxcxKo42Em1MxDxeb02Fv8588oOz8TuOjej2JnKhKaIAqD42DswylfGFMs7kEdmkftyRg
y9TSslouvSSHNX1XL9aRqEu81XeWZNgxpqwJKP5+FrlAbsn193BhZLPygFCG/vW7XvZ35syunwW7
qBnj48ZsaFNDAbuS3g5xrHUU6qqR1Tj9pvY6EIvl35UwsEUjJBTAqpQCaYkYkgmrlhrPhC8h5024
MqYM6T3yE+hpwDYZXr7r3pNpKONo+vn2oo8LlgKu9sltUpe99tat/4PP8ywxHh04baIZ8LHC4u5D
g0yETowr0t8sQdNsYbTCOt5f0LmSGsjef0GkcNvIvTNneEB3teWZHjRzqu+l+WxuDnt97MHAqLey
8QdnSUZKjTMqsH1NiGAKaUhCH/wynhlvnY/CobbdFI/z5GMxAmx4ZkBRTOFULRkajChuI3WxNf/0
UFd8lhwGvDVMrmGJwbQ7dXNULp4xmHzaLrC78M7FWmBai2wl5Pe7eSSrRtEm7zHRUTvYG3O3M6iE
+lT6Bu7ziBk3Cqb7rN+jNR14FWOenj/94iOUEDWUlmVNDa6vta4Y5kM7ycGFKDx/K6IKaPv7pPTJ
V8jGUXfCMtF+yGY6NKlJ21h2Xd2HGLXHVai9kQZQtrS2v6jVSbX8j0EsazAg2d3W89OSBIYp/Spb
OHLiXXXrIgPB8MkSRfvbXF6OBJO5C1eQtgahioYdUl0uop3yAqcEqcZ51U6F0K38WvOSpbDKu+MZ
C40TYfxlGj4+acf4eOMlmgnpl+mbGYfuA/1/K136AVJzpRjQ5zA5HKRjLUniPg2uMSY5gYasOX2D
k6vE6C9lexRINLlFsOf4Ukgy3u2114/btB1rjKOEQdX/KzrTAGLu4fDx6i0wiUqBaVmmaRygWRPZ
3+2exSqXt4DkEjzDoZnzuXo5IqZOmHlxiCLE72JaPxZ8RWg0zUGKlXXrM2aBA+290QfXQGhiwgaQ
YkRywsEUFqcPWdR6tRAuXcJx81zxMhaNaaJAay3z/PprJNmOzjVAHB3ChV0InglV0b/INjISkZJD
4i8+fCz9CMm4oxdzeAMWG33/rqSTG9nRDWsaxBSvGLRjJ6rdWNLVKCQ5+F2A7T/kETqCTtahjmfE
kmlHn/RfphhY9GimfsMNOUX1bBh4pcKa3SUZ4RL7r9IMc5eAs01FfYOSwuzRMpsCX/QG2kLhhluN
okCByyh70LITqPuAJnOhEkMTWGogZhTanb7EjiqKe8KeyCygeZOOt+4vaiA6vSbLhhNciuZLcMjW
HMRQVmrl/XPqpTB6OD+0DjmPq6GV4Ie3SAi6t8jClOweKTDHYBNbr/uAuHCU+G6/F+k2RutxkggS
LbRGre0rEzuaB9M/i/wSIGw44VQZtsjYHy111VpsvhZJ3+pcM0utfIgS2A0kY4YsVbInTSNV8Y7R
YRdLffEOfss42MiXyw9TuvI8u2BmSK7cdvXGl/nWBv33zU80VlYigGWQpTv0e5yHqEZxQ9acf0x/
1dCQ6hDF06dYY53oBqEkmu3Z/4oUjUomrKGKT7f3V+3iY9ZNQE9HSblhDrJgBVVN+EO6rRvn4Ep7
pf3mVyd5y4XrCs4/19QpFdiCL5ayMQOLHCpXzxvppdcJJt/H0aMO2AdBxGxTQiNrmJvdZsDNbjBH
sTNBQ6MUKjkv9GUwhb7QwNUYTh6TKnn/japj9qCW5R+OpYhgLubd5908gTOEqyvYLuA4uIxd0X1B
Uo2ayqwCFcMubytqUzxJWGN/Lj3G40HDiSa0mdgljhfkBViaHXlN9kc79D2SxBarAsclFHqh1tA1
wUMFc2bfVkMaPKBruQv0L6ExZv/dwuCjhcExoDVBV0Rpm0j81tFp9WY33orn4if2C7Q4xNAxa7WH
P7toDRLh+Ah1UeoVvId5B77yvjzUs8z4KnaEDXwmBVtaUMA7CumM9hdRMCzjhJLjZg6zrhhYdL9k
V2TM4tZjZyV0mf5x5bX/DEAo0GdgN8WBA6aH6JrR+CLBRXXMQhljOZOzegsJY6uoaC7wHM3QMf2S
AabfPmDOhgvqYAhJgu2eEcgvv8VXi0O4nyHPS3sICtyDEuSVPfqqa+VVx0+cSKDUuhxOXuk7/iAm
Y9+i/tY0JO3mEjojzyWufa5xRwawUf6jRdNx8im6HVXOVZdRnPQueMwSij55pyKx/A73NuMEWckX
84LwXtS6BR/vFDye+nnU32E/8SxyTsLjbzfRTk/QGUNUqTlZQ0bZwQP9Po0SnKtkdDps9KSo12lS
adLvKVcI6S5BmVb/PrH3X7C1+d720XSCbH4HUhPE0xn2ILN8hurzcX86nlx7234ACiarq9nesu2z
DLr5svMQftMctBRgws/0Nb2oL0YeI947Z3btBeJ5RUyGdNiwfkuTzEPybky/2GlO6g9byimi0DhQ
kqXRHSTWTkn0A1+KOt+jr6gKs9gwT1fCdgxS5Yo+vFuYEonzv+1E9LLtNHJWX3ucP6GsCVsGZrm2
ciJPk9NI9SvE1v9w4tik4iityWnvspyRxNvFWlqjnK+hi3t5oJJ6Nmrk9n5D40SyQBdmlv1HcpBT
DjihxaWCNdLyrjpsAZ2y/Jx9E5il0/2cPa2B/UljjfrZwpJly8U+AOC+8+DH39aCN+g3FiuYg8LI
TY/TnNki25O2k8ZNJ7dFoxsspHH10ugdusc6Bnyrjxuy39sStcfHFerlq1TxTF9ejQHkdRwcTYiW
JBxws45iNhc79I9ABAA7TgBNK38m8B/AuXhebJbpB0t191B/hGDn6PUzx8dVOUJByjvYqrhEpCbN
+kfqBz73eTeOa3r8DxCHkDIz3xuFQNt4TDgrsk4fr709MEnWukbSlirkFK0bed7Ie21P3msIuIJp
LtP71rJch+9W2t5ryZDu+ujGGVsU8fh+aWmEwWbkrNW3/oVQXjF0D7cQ/tlon6wbijDizTS3DJVH
BW+BKW7meGN7t1dpLVGeK+3/dQboTyG8/rOLzxUCDIWG5+G+9AUBSfkU8g4K9ymZ3Z8bloJus7CA
XfPeOyg8jjUCce/aSiSVORRI6sPJi0Rcm2FgGCnij1od8MqTSyYgfqMeeHxvhsIXA+8RKJP5KJ/E
DQDMDyGHvtDIxJabGQG2rfnEOWr9rUMVjFRi4KngUrSFkCx8laexw4QnyKcmNqd1RQABNcEHf/J3
jwQ+NlsIqhOMYzu3JD/doD/7+qBOjKdiYp2RU4gnJ8szSuRda3fohAJilLJ9koyzrKWqrfDUt9KF
sy/FsiK07O03/wYEcx59+kgB4wAPHJpx8U6FtbB7X8wVc1SKaUGU4ZJC8mMj691wLKraLi+WDjUU
M8uKISrACV0R/caWvJPBlegTS759Pt2n4XIKF+XA5SFFBPRgG9LmyQf2UPRxVfRW0fUE0iKJDXvp
GcPQbfehCzzIXgF5EtQ6sPlU+/cDDBqYg9hsN5cRRVTuxQAX4nLz+uiDiEvAXzBvOM/H98++1zSl
RHBEg0tAny9BBV3I7dx/LMjer16o8ckptk+kbpmb5+IkVZdf1dOZ6SpJ9nmNFbObzfny3Akw0XyZ
vvu0CFaNxhgqCFzIyM8WnLt/RXhN1em27pqw4I8a9tpqxoPy/deiAWg9/c3sMaM3NRj3ZL861nL+
fhwKzEMGEBLLX+oGFAxb5XkxwyfP7T5pxUrQWwp72BV54zJihzoU1jb7uzbVKgsc07jcccq362sy
7c+4XWM+H4SFlzeNL3x5/wJwGQRUyJ56Rrs/IAqLPeLgusCCp0gUqL1X/NmhUSIEHBYTjhRIOBfx
HAfdQbgRPDh55g08qZqMyrHuCtenoW+zNGSHW58XGJjFDz7o+bAYTNwFWlG/hUwB5GYLgKNakBU8
qdDo+uQok5s8L83djKFLNvjE9tEMEUbBxvUJkO/xm4nt4jFautjqpsRVRmdQ1kubwi0V473mQ8pT
ViMr8pKRwcDomByPntww4OjqD4cY91CYwlpDdFMMlnhGRJnHc+6Gju5N49B1fKtB9BoFS66zfzq/
iHI0jL6+nNKywIEbDdn9Kr4gY1dHqPLJ9c3mllNOHg/zoPpV3Vb0A6xAacEb8IA9JeZYNBPSjl8b
xp2+CnQn4B2Qt6XIzEzhBcu9GfvGFkjBXHheFePNwAh56v9GMZOT2rFxyJSW3epQhVxg2p3kp33A
JBMjL3UQcTD8mj88MOXSiQ3nI+wwZRC98Tgwng5EN9oSpspABQZ7Hww9J4qXrrZLl05uNI9iVUrl
mHC2KuCUBC7zZE5EYq4z+CdQBURBh4GPpunRnG7YD9+PQ1+2jNhUcGWxqMajzTBLxPB4LA1Pnj3Z
MuDauTT5yOmGOCpdQJZjCsloCEydLr0sOvEtVVYOSRwXuqaH3sHyDoe+HkLtvsWVV5Lbh/g3HLBw
FwQ1MiovLT8mFg0ZNjMvTNWxPpSLd/UdhF4GnDOAJzqt2/PUSmBuZkpexWCnVttvhkx6Nqiz741e
C2oZGuELyxIoWIesZ9zXi1PQn3ZgsFsBR8azxKTufY3UsVRF8T9E1Vq1k+FysWWXSu4kqMZvlqNN
XsKbMjesSHh4HuA0sAurxNjZnBer02+9bE60J75W5g+QSKogYqn0fP9TU/eggi0phtH/E80tpsTD
+n+xKJOh/J3wQNJQ7UOQ/CGI0hR1HiiCDYMrbpQ8yJlmsvsen3nsDrPzD4p9wgOapT+rc4aEp+X3
e1yBHM3HzyhRE8ceBsn9zylTTnD+XYm0vlyn27T2FzCOuL6Zo+GmZs0PngOZR+9rjWkShzgEY2Uz
J+X807HYjUa77JhL2HkRygjdLXRC7dtP9nW+3wKYZPFo5LTwcMW1w8oCNDL26m8zwnZdCqVI/mg1
OIwS3nOWLGG/H34zBoZQtveHwGTQGdGhe4zlf32avZwq6htWKFn6cZffsjPKb7ro+a37/vKZpwhs
Ufqazb8LCmM+8cbwtlaJ5fxImK7ziJQedzPyHdaVCZ4c3KkN3QV9wX03NbyIY/GQzoHNL766lw3q
bxz12oYsdeVnUg3NRrw9P0ta+OlYez4U9WxSjILNNAptp9QTq7mhGSFsBrh/NVJMd/a5h2I47jx+
nQ5c/koXcm/wZD+zgReJU1GkSQnrssGNwUtrnn3ggKcZTDCu1BzM+tXzi2//rsI1tWyDH/03pyBw
f4M20GWx4UjkVneRGw3WF8WvHSsKU/+B03SwZQbVTA15eVRFfUkHMQArC9dBaFSwxHWgZmMzHz3c
TrXbNcKRSGKgp2Go669CHh11HGw62k2k9iNV3ZzR95IPppKZ+hs0kb2RJGxSioAA5sraWpHc1KNJ
rmJCkPReBWuQjr8VEC79xbrO93/bEkqOzIVlAnKUZqTbWRjqZFJFOiwF/6EfIT6TSqWVQfFkVmIb
x5v4zbC3OJ58y2GQZx/oZzBB3GnG+zKCxsGk0DvyTAv6YW+wWuOscI/g7K7gq2UO3sUe0gqGDmBD
uuWC9Wuv9dntd44AU0zRj6H7knVsfdw7kxOr9taT3pKBeS/6zrrT2PqnRN5YPj1zNEpEatvuPXhJ
oiulrKJhD58RDKAkMP/kRt7s6cGscUJV3O5BusThzsp2iipA7wXONAovR/vYggFGy4DE49817RBt
6OXeCDTT0ZRhECQftxQhRfFf5TDw4eVor3XpVIetI2jXeA0Tf5Vfswp4ZxWVmL6Mx0nNWOL9ua9K
85uH4gLEgKyHJbD53OXhSTQ18qGX4HVpuM1opb1Dtal9pZBY94w9NFB+MrtK3GFXKw8UQX0Hl4Ul
EKAXA2LhzlNHP9p+0GHeTPs9TkejkjMuygXKFAomMkgH1dtmj0cdb+YMqNUsoNcoWv2+nGwRwbux
IhTqYeGpk/N2M1twvI581PTWWp+ZYoG4YUieJju9X4xMxgPHRCajcjTDB8AuiaTJFWc1WmObbX0k
0hvJHFn5ddbBGDEgiQccM5vFfw0a9sh5v3rZmdwsVrLOvnXy6woBPwD+HPxKmF2z+wlW2wsjteca
mGuWnX57CpWmfj6ohaQLW08L/PCOFGmtOeajWr9iH3SywhwDBTCADoyTbVLLqEoBcw1DVR0la8+4
oYytU1metMlUVl2r9AfDuahHqcscKMeYcT2l8d/bAWTxPsbo9xORP+NlhXtnaGXwodeWTwBl2BKS
G/kukMh/GVm/Di3v/OJStp6puCH2aAXhUlPt4uPpjdtc5EWcrzLQaguTdRHCZm1v9y1HdUtPZyax
1gJoj2eO6ufZgFRGcckFOag2TEQBTfAVChjk0S8M1LEDdrp56FQkz8hQSwXpJKxjkhCAKRoQPGI9
r5PfsbqmZoiQutD6fcvoZVK8lfB+7CzdC8l8D4c5h44dwKQIEPgnLEux8w7m4zJSdi4NUGLHQDKw
g5T8eyEl1ku7P2A8Ngdz08cpCMPv2pNIOrj4xiylHMdZ944gubRkQCvrxsLOJmurKUPBkWovaglr
crO9a43Lnfj+vEYdnDCw5aAXtj1Qs7h2tidSZJGsyVv1K1+TOYGSYUCBupsxVmkWBCamrth5Hq6D
IviPHjM8Zq1z3Vurdugo1k3ysVX8tid2Nmmzs8uPlRGALJQXi3DnjGridT6drnHHmnzBQZN78NzX
oPNVRJw8R6qlgJkl/s5+CMI7N7pELjIWrj1OsdoDjpi37EqTAEngj/mbbw6pJ2TANFfd7JF75tm4
nnchBW14/+wC1pVGKZierVbuSU+6PmMdkp2hl5DTw285JX2zCm/nSXItiqDqBlaD4/ujKBQ5gBD4
WGH73WoTKYWl/LMOe8Z405A0EtqZfq2hE40SCjzx9xgO7+JO84GLx9BEhOtFoiubHG23zDX9LFl2
I2n4BesFToq6xjF6OSwHv2/nxRS4OAW23coSnY/OrGQOltQMAaUUYPKWo93HzLnNkiUzisfoFGoX
ACrNFTAKGTqd+1TIWjfw39PeXHXV21G1gJdkejkR/uwy4ZzCXmrEobhcKYmC5Vnr5LyID3xIAMAo
XBBOWD4rK34POMLQ+HHuRWZEmkS1pgOf97e07fGwAyy13xLRU62gbST7yu+N0Ya5O86pOoP4mqnF
UkOY9pjYQtaNH2Dlb8AMkO5s19PYN0D7PijPCG/SUgGJs3baPgW5kXXdfaIgX1AtvkYOErVXi0ZF
Sg+IQuo4Up1Eq9GRNPriZjIsfjPc2NX9ksV1sgzfHKVF7gSVB5ZjYZwBWv6fYpOiiOEBANKvVtYC
OziKvXlSG9/TnzIbkr6+2xU+jUlLhpNgVyuxhZrTsRM5ZrXQUpBdfPQ6Latz0h6UQHH9tDNpAbtv
i7yAFIozKTgwcjzZqfqICX/Lopj1cw97LpsLkpEI2wJfvn9l3YBLb9tD6fQsv9463A/tU7R1x+Kg
efYLGdAGgi/3CH8qJ0tP6+vjgXFAsCSa7hm5aOo2XvmSuKeI369ad1xFQa1aO20VNC+YuepiU40T
LE6Fgr4vdqohRUVVtdfy/mzxYOvvRkqjf0FjoU5UhPeuE4PYSCmdQP3Kb2Jq81PYIMSOxIZ44tM4
FWk+CJnpalhe9AsQOXVkZxeybVu27dKuLnNJq1U8MCD2uN8NvZROf1CwDrutZnQO8qgiiIzlaQNv
4ARNVB/1l1WWG2dbzbpvq7K7S+GnyZi4o/ftQstw0MS6SpF/M0caeLL64wpNUCOJSTstlnaa5hEC
FyKDGGsDBBWm2J8yE9QlWU6DB9G/M0nIsWj2hXonL2d87WcI7Z/ibOefmfKV5aYQiw1g95yX97Bk
Qm+x/V7n9kq9ykMqmNHFBv1z6tuaBrCJdMcru44XbZkYYmtKMzWG7fYrmKl0dOCUeN1p9GyAf5NL
kma31+a42wZ3s6jSJi3rfzo9/f+dPqMSsQJQ0wwf0PyJh0rBP6t9AC1P8xHlFJ9rajQJf04Esr+Q
fCmBSJmRVuusdU9yT0a/Nc/chcMnCiF4Ia4wRTIIadqNF0rQGibdc4Kgx8woclr4FbLnrYL2p67k
I74No5lZEPIxbIYFNsfN6CU3c3I8a5eCoeDHdfaOsfFFujMiG9ygDINlWFWV1+sEyQ7t1ACIoCgd
l0XWICgoHVGtKDXNNQgurV2dWB4b1XRDuXdliCACnz6jRBlGOm96fQ9VN1Zw032zMozP1ol5yLgH
SiNODqqAOnTcANsZtZ8/XJM+6f/0XvYA1iy0I5G2KxBci6UDz3KJ9OQ6KVg6xnau0dzYXdxpa7uo
ABSiXyP4qW7Zfz4YWpQUehAP3wvVaTgo8e5gE0AIZ/cE1BnCk9+1Yqh0L5cnQ2dsJVDsC01Rlx+8
KCVZ8YVxmk2W9AQTnZZjEMFgPFengmIwVa6rnOViLQenqEznAnAZSuNd13OslDtw+66ZItSHPzmk
9vdXQKy1lhdHZloJkkTslC7I79P2sQi2eKN5L3UOhqYkf7dYzQtoRy8oa+FB6bR30qwyXcTDfjNC
axHQJeYA9YkEOdvOF21b757cUugd3Mgc11o5ICteBN6+cpvEFSvMCuK6wBTLmc5/aDB+bi/IUWg8
d9U2ROcJpqjN1bmiEgmFHshntMo8H5IgUEO+tPAtIpDLRGUmPbGUqdQyAie7qleoThn70/OHPGZA
BYbUu/0qpJoKLanPlpDL1n4/OcF7ZyIyGIHAtmsg2t+Ohu8r/vYJdUcAvDgiOLGKEql4LEjQylZB
5kAPC4uvAxwB4oCYuLIB7kmJuithEhYOXbGeRABEcjlRMKJzdpau1I6EpoENYtXTg3ghUQHbJ4Qx
d5bs4cN6bXWDpuGZcBYh0H/hJo02g954a6TcTTlGjY7RS4UbIIFkrtEyQOddIl2ClZHrnIfpbGhj
kTvN6PUUwFSBmVUvrW5vcW1ETMW5P4tb0R27UJ2aQgqnOWtzMpW5E6JTPnedcwtUo8FdcAz2Jp8U
W2jifhCsifrgQBB3tpLDADYxSYVAuLHntFThPKiVP50fG5yWsGFkrbdwkSoPcF5v8098psN5o7ab
bptqBCnLt3TKdHCGwPKGCraUpVtHjiIl75PhCoqDvlh2b3qJJ3Xn+KJFqJQhHf4w4R6qG6TfL7gA
BIwZwMcW87jGkvbvWj8jG6Dulo5ZsBB6w7bLJXB8/+dpPqTIPGPBZ01hl4iyE8pSK4MUcUr0pQkx
q9F7hM+c8K6ltHebNDhHnqvUwynACbOxjsMm4CT+IG9s7WQRO2R7rv607IRqqXHI/Xaw8RSOduMO
wF/gvJG0ANXFR1CAVP0gB529x6RSIJe9GEkCd/yPCGSH+DaWbkNjGB9dwNayYKC7rid/6G9ahh+e
BB52idjFM1GmA41/qlVb7w7l92ZZ5X8n4owHfnUIcD9UOrUN7p5EFj+nPXWVz84dVis+ngV05zgz
Nii6eagwUSmbBP432bFI8cRJO91IJdt09k0AEYRTxnSKv4rxR6ug0lDpdpJ9UsegppcU4NsPlpWR
w2LBomt/NdXGnPFg4tHNhORqQAt6UF5OxR1zboSxkTm6ognNjqiAxNpCXS408FsmQZghrE92BARw
Z3t+mLiR/epcDbaGQ6p9eybO1O2UsHC36dBN0h2DsAlN9vmlrk6XQobHFI9EYJn7HPji5CiF/7Nt
FCd6O+UpYVwiFFbH/icOOPrALKxFhkq5OHcHXm3bNJlRjDfafSvY7tCuAu8wV5N7k0MN2zN0AkAj
GgW1KJ9YrrKkRUpTlxFOfX3xM1j+3lPxkwW1llycvshxlWCpyEejlkDy06dpYPl5phmZ4Z2Rwdxh
rGRwZUOh457S6FBdEJmYhUo+ooBYntY+IEGMVUZZrS4M0TqtDOISCKqSnSLOa5nIrdNjy4B6cxPv
G/5ZmZhWDI8JhdEo3BouEMV9i8ODcrq4SPUeAkikC1cbL7xmgqLBBzNxrWQIcRPK4b9vRW4yShHT
+x4u1X8Xg5zuBGTwzVJ95BZcV+guUeAhleasHreQCAuR2Etqpo16vZRHpRZF5b6cd5N3HHuGv/ZL
NvejKM4a6oUq+amJbMEEAmWtMSJVESKfbsUeMIzViJf8/VYZ3VF0ZfYTB9es8r7X5arDtO8ywmkZ
CjVy09rOcR5QsQl/W3Dp29nidfE9ZF6SORUIJIRBuQTGBe6miNPu4ZtZhTeaKbQUtx/gkmHS/VTU
gavYScEJQ+XE7NC/1y9rKX2kXZdbO/s8Uoj/HQ5v66KZG+gOib2vRbEdf61oAHBIYeix802wrffP
SPKHwD1QC6Ori/8whvA+xMmuc/KoUh+0s+InqCwNdUDGVmGFw1KacohKbiivai4SdZ0v7rCp0rtJ
ribanztMHRDx2BN6BRR5n26xU3blhTN0NV/tnzB25DQ9LhVTCXeiwuoZASPjf7SY+NSnMQoJiyuu
NlOkUBUTxH9YGe5NdibwTRqg2oW9nMer+1O+MJSeyt20n2djc0PTNRY019tR/nRyPjjV+fmWQIV/
V3jKOJ1kyovGheND5ovTr1FYHDzcyBQAn9I42ZvhivsW+CEdLPMAZYE/I1bXlL9PqMQhcYkuThN/
nPF4G+fngxTW9MLQJeSAZ3KF89ge2xwlLKWso5EYVTjaroFaMwrwguHoeS1d/K0Yeb2m3Q0eJNCq
nlsjNktr3cIqhhGEXSPAGJaxizh+deR0Ye/qD1Ai7ybnCiDLUx0sXnpeNdq5gvkt+lONJSXe9t1D
Zn+ECSTagpMqHz3zGzoOCpUvlp7ovYiiwF0My4Ygrm1+mrLlgjbOQYa76RIZ+Y4omLaRd0T1tm79
kpQWMYYJ3Lh3IK0esgm3C4KB4LGagzVKPJg83BR++1zhcLaxhvZY4jZnDrdvGlGCwKFNy6ZnryV2
ih/+9vwIYJFLzoSeJOOetH6Wh+IqQraoOqOV3furQG8ohkBzUU9ozavw2FyjCRgZ6RTvOh69OpU0
3X+6Fu7spB4v4bIo/0oY1vjfJ8XejkpydyoDj1m3uTzo87q5XHt/Nqp48rQG1Xy1fas54TVckdC7
AEEPeGTSrHsjkzZ0/E7p3DjV/O4AbOX2TbkMBE+7chjda6nz026eTW6TfR1Oktdo/v91kcX4+/65
76AJk/53hPibOMtPpn4YSyDctgg/0Tc7EdK9fUglocggkyHXz+k9xk2OT8qHYs9OcZ/vyWzqt4GN
sZXmse10KlwdQZPvT9hudOLrets1oj+Fryesz8jg4b+8wXBCimvDg11IpFhxsJ3x0tPTrR7BwQSf
W+QBKp4pokPv8guHWSgnxgZ19Qx0m6LUPa8jhhPsoKHpW3gF2WgNYeXW0jy06ejCCaAUkSFc/fD4
6FB1dP3F5JXqr1CCfz+CctP0Yjeesb1N/hkfLRyIpdM/yaKJ4AcA1kiuCUzOHlEp7T/UOPE7ZxTb
ZZhOvIRL+70zkTKE1fYAZ+mXw8T4mKVpurKpTkegyeAFldtiRGsIK+AwfBZOn9VKy+dLlcDRZh5F
vrfgLhTcR/hNakZdSfti3jZf7AnHcOqOAxd1SrUHpfe2JP7Gd8v8OYKM5bcWTOFKrrn5BJzQIKZp
zwKKMunB5Xp2j1MXGitnNNbjHVrxos3oYNmfr/APmwNCn2q1EHM/Hj3JU9b40gJQu0yu3cb6cBNO
CEq/uKKo6Mmjo6MPjKqDwdYljVZIkZfq+AC2GoI9Iau6Ow9PLxyP50Jrlxt6I8VUFWu018tj7yWZ
0ramVskBy5RONEj7Ut8ZxUHDdthyV153zgBzQGiziBmc/flzE7YSnFqiBmLo/mYalyEpAmeMp30i
k0viAV9HoROjVnbJNHNWXFxe2LrrLvMTjDkkJtWBfgCPEYeubdtCc/hiwEwo2aMGdHbomyjke1h+
8Ee4QiJVxtHPg9DrlIqKcxOco0l9xegPTpTeIHD+KLv90Pv9oSRMQkqshWxrg89+zOpIuu5pzmNJ
EsahyelsA6smtCzugplqea7qcTKQEclbrLKakvsZIoK9vi9jMdQhoH3TcsPrOb8J4beLkoSbgP5y
9RdjA7uBa6+SQqzJ2ox7RN6xc2IEojZSC3nQV8LDpDVxywOy8tXaRGIiCHoBedgVLubiga39YUCQ
NT0q0R3H6+vKA1m3H+s5V5NmMzpxa9Fb50ZRq+i97II3r3lppki6ioAfugvM3ZtxOnbzIduTurkU
UQ0Vl0ue3gpkoODGSATHchHwNfi5+Re4X6FiqeE4HEDh3D/N4VwQs+6G4YrL/7x+HtIiOkEjcLcI
kGYcLI/VCF9dnhVMXuQloRvqomwZZ4TZHP96QMzrM7tV1/q/2xxYthFmGvn0dIQV8tULrqvl61Pm
RmlIzXD0hGCf8xuq8tMOadENgLrcPPVHUcMs5qAQlMdthJMxThts5/IcGVPFSmb6ldqKyd8FoyAm
/30sgJYyhNyVb8JS6/U9IxSKvQbNm2eRuHcnqCggzWNj05gz1KRpg/Q9YIT1p3HYpK8rju2ik21x
pgOVDkmHtdV7BkaM47hqilYnTHRuUeou++LfZoZIO7fcUyzMU2F6NzUb3aFu2tFaYWrrAv2s+kSr
BxlQPzQ8Pd8vRGwGXrXSelcgx+68y9fPycUunwhvCSHhnULHruO5OxKuBHkzgZWDVTHKOCCR6woI
HXCQYcky3sEH2vQKY3ueqYwOaeLCt44a6beMN+2AD2TDLBQD3ktDDt1InHZsU7HXjkFCTintNBWV
Nm7Y+xGakZDC8ags5BWhaOQM6kwgrfFtACN+8bBPPmnbU0oFyCyH2cGGaWq1C2LlEOK4uVGQjqRN
Apu/Czk59XOmxpuSxqi6eAkpu7OjMYlSgM0EBu9PAFfejen3WZOXrvqPC8uUNdDlbYGS2NQ+yfeT
FUA/SwL8EmOeFt43ylQc+auvS8pIhiEvXP2p9rWA9piwe25mmooA94CLugwyjKNLfmQvUeDsFfTO
NC5KZQoH7H3dUDMwYBjYAn/qogFWe4IqUApUXe+9xWUlvtLsdJfnD3v1DKTjY4iyFRu/wE0aieSW
dC1mOrKx7cvBnXt+cw2sIIJ/2O864Ghnu3tQDAIeMlD1gymIGTdJtvgxGPGPklGmU3micU+jXPDh
w2iCMYpR+e/IQzJsGiQHrDslk7K0MZlwRJz6CCq/Hld3Ja3d8UxTMQvz073a66JhhkM48GTPzXOL
IZ/7onoGujchWnKZ8BbXqA/a5EipcwIU5J1rAhEncTAPKWuzAIh+79F1eZI0gY9WniHaSy1cWkBh
7/jCpfjgYOlu+ZyyfjKGRxph79LsQuQ9y8NfJK54mMQwBolpZDbfVJA8F9NJXGmExbazdXojvrkh
imx0IkOF1zVwj0p6wm3D0aw0qIJmhiyaJbpHluu+SwnUcbPHyNhhD+uE/uPtgndppS1B/pZUMrBC
gHQrFB/yM2WgyRPUL1YmHxAJghUFc01pvtsMxAkCa6/uwAEQzN3/dKQmVB7k1Bkq3BwB0cInYgCJ
qMeGnHd5lGyK/d2I9vZwW45yl7Jb9cKiIqNc2RAU1as5J3PgSE0T9K81GvJ0TLR5WwFFifAMcNcL
9xlGpNazxJZ6TagGzkE0nCJFBPBBIeA/i45ef/6CgtujkiI4jgLzoidbFdB4yn8ckMtmQqwAAeNK
/dCPVnAAacJ3SmIQGmhDl1vW055mJoJnbir6UFCyAdxIAyDvqysgkI/rqOFiqWPlwfsBc60kDxSl
R7R7IBLrHHRGeZc98mYFsWU1cbJngiSGjqP8Y+Zjkn2OCwVRc8jgycaHPZPf+Azd615ray8tQ9rT
hnvSi8r1E+9mFZzens63Wn3cjTYj3wRaZGxHOFh33eMiuL5nH93jF1hZLsEFDWFJUOtJNW4PkhlT
iIQTjEtfUbmgmLj8NUbaoN2+EAO2hURo2FIDcOpH3eLP0QDi7Af/SA9Fh3bULJcgQ4RB9nqIMyIc
BMldfOL1wHSAJRZc3tRAraBK22TE0v4i0nx72fgMlYXUJhKg7I+xdUVAdcB25AMvYzgidhQM46Ap
6qMgOkOkJ5Hoyb2m668+FMCnEyiJMu5TznP4apOGQu+k0skjt5pdi94NxYhKEKL6aOsVotL9WIwU
2vfDFeK9b+tIx/mLCMwfU3cF/Z6wh8LopS416N8BAzZzDFMvoSoxezMDQaGzWgsdjr1UEX63cEiV
sP7KyBGljATW09d7cnYXt1ei7v+oSBMks4MWbuX29jrFkrxj0i8HReum3WDLoxhbrFtt5gp1uvB+
QrQyyUjI6BjJPvHRm7Ezb/mwz1dvRtMOOVLp6GX9HQNMG5TSQVpZ05o41/sPu2KhRLGaOAJ2RR8r
Xr/TQqviCSWp86w0n+6XlBq8vFfG/eymHymRUz9xvPQugfVq48vCd7+135rFDOfBTW0krjD+WeYd
Hu0BaYXREHE9lKa4juPnxWh56qexNrELjtT2ncUHzqBc3DkAkh3z1Ng2OjACMMnLIRkPSfG293Ax
RXmelf51Wz8tmZFc9iR6+w5yX0eNcCt4Zi7YWEW/zRg4HK5NB7KJPYT6PEg5R0a+5F4/DePHcdAk
Vik+bEssdbX2rY/ycAwfk3x07ppptAtC/H7VQD2dqhQm6yvKhQhVSWWU2uI+ZVpxnxp+UQkK5PNS
1wv6H7tYSE66Z7nSODQ01AUkkkXJmJx6PPgeWDwgAqtZOrwcjx1g43dWBjUR37OPFuX56slXrtLu
TnkKVtiKb6Kzz8kEgruVHvvk5E3wlyz7IguNZhyWiLd9PWzFhmY7zGOjtGWH/9u1YytyrJgu8MwO
bzJPQzvKYtVCiVZX6WVD5NCgPsjD2bCGpmN1MLoBrhSBt6w/x6ASZUXZGPzUePmDBk8F9cC+1zAz
mgKOWDirc+OK1xJYhdiUbcDaq3ArrijWf0qTxBJTGi/nFCsqj9JFdMwZNZn/Iv3BsZmUddSmGgR3
1v162Vbenhp2M9bt2WuhFGRZCYCRbCdC51vnRtIWWLy9HGEBHQKdPOfs0fyAnPNt2sGj6dyfg67o
4ZxKw9iflbw6yi0ALWuFm5KftYCgtCuU29tKEkTwJ+lsjyOwZ+tq8JvYwOXMs2g527/30vFuxwT2
k1irOMOv0b2IEAQo6JJ3hBcOOTQbjQfHUHZEWdTgPTFHzqbZDO/bIKSeV6QypDakgA7MZMMeLiNj
HlZQJtGODZGlPj+5j8GpElhtWH5djHvR8Bez5PyoHG0Y0B3qdWCgGHf2GWNwG6AVTjnOpl/oydyi
o0pidqlqRaViswN1UsUvKj7O3s0uHJipF6DYeX4Exp6cvz4DtZ9A6MSXPvhFckmAGscGs0y/W/Xj
9+J7wg5Q0enEbef6pju06pxWdngk8o3BN0A/A/6lD2bXFQF5q8HaJ1bEthpm3w2spaJQUpLgFrmP
qw9y/f8YXlqoKKHXajTiU3pOFC3WAjST0TmO+jBcef3s0tFypwsztnYeOyxOrX6/mk3acYLB1kNA
3C7vY31HLTO6O2yI2/FFcKsG8qByqGplic3cnEz+D6OXlC74uK7olUHt/G3StYHioPRrs3ipQ6aG
05siLkZZO2bX0ZB+eXNTXYzip8iO3sUzFMHX6m6tmLQKx1EVoyXledlce7Wm3lxZ2guixXlpTHwK
uPKr4Gf2cjdsgG6PLzwC+WVI9PzZe5gTi7Y2XXnOXdjlPTODVQRV5nZ0LtZbLyipPDSQ+YQjtdf+
t8QTHz6Qb2hYFaHF8/Wk5U8qYxO9AY1wojop5R3UVlsZv/0z6qcPaCzr585CdEJxPTfEVc/uA6hG
VDJVIpjLP/8y0/Jgn7k8CNmr9VfSIEzqfi6xtv/xbSo4P35MXXQ+OuKNyfLel3HvVqk2BBIStQzq
CYTKFyNp+oNTwxT6/rv8+zOagXtMfVyCahP53aH4vRM47xFV3AptZzY5jTT+xkJOXh5ibaGHFHeo
ykbABXuff962Q+6rtDT8WPy+JWtDLRMSZbZblr3/vEvTNHiYrSgeDM3PCCM4ldFCtpIhvxowWvJW
lG5fmQOWPENsffvyHMHfkf1IsP1tdh6tQ6zGMz/8uIvcM8j3lYhjSJJg/jWw0GZ4Tf3wCzYOiWxk
iCxsHbkuE87aeecwMMMpDFZVcrrC3Sdt4URI5VRLwb8zs539CXpUYhI+A78iZpAO7W6/TV06lHuh
IjuDMlF1kyE5o/6pK15sf8cqTL9KjtFaAXWpgdWrRZnoPkWc5Fnaf5210L2f0PJtujRZu+TYFAEg
V3e3xeO7LE4zNPMPEfcSBfr/fO4aqDMASxaDWC4L8/aYjfyO5neTxJk2rQuSw5ne+RLczDcfcJbv
JkID/uSapNlIBhhFof96YdXzN3ehpVZBMQXVr+y1yR/n3YvUpzeebO/ga3/4326dfhWSlXqQJ0D1
xeBUBoRkP8qrWtoN4i3X+4fp1NkNJBJcmtf1lPwOQsSTKL6pNVaAIBzxq1lkP9E6uyxt9alj3hgQ
Y4zaULxVSRHHlwutgnE7BqS6EPHG3gHsulbk9QCBTiO7u/E7uBgRpke7C1uYkBS/VZPXGbvY0v7b
EcouWD5gUTFrNYm3OnIa7N2Wkp9sW4MPXBYintsyUvMh3OH/fAEaKMaKKrKw1F88PV0ouoVfC17+
nGkMjMOsvUr/O20MFd/mWQEpYWhvCUvJEmq44kkpCV6HiBmaIHlCb3oeEJO+zjnjG52UhoMB8Dzd
ynVF7Qsoj+ZOxYktJBpwxIavmcckUqO38vQLXR5lDKWa2KCkfb0grifjDOZ2HjVAx9hgfXhaMjJ3
X4gLWz9wSOkEOwDi3hy038Soc3hoAyoJcuBv+1U8r9vkknRebvuaymZUQ35zdL5aCCoz3m4Y/Rdo
+0aoTbG+ItofW0cexnfh1POgv/L3/PJhZOUbAot5WrUbedU0SI7o9jmVEKNvX95uW+6f9U5Bnv4N
UzUCNGV+mqQrZA/fgcYkHzgsHdqUbuU5YqvO4lN3D1R32Jf1dm5r3J9W0NFFU/kEZH6RNnrQGi6c
iPfK8ocBWya3NU7hI264nZrfMdR4en/cHxeRLs8YmdTOBElQAwOqA78UkzgxgjLYZ23MHgFatX8Z
VtHOWCsZ8q0Icb7ZExSWW8H27TolneI46fYFK7P/GBjsH7QMVLRQnrqx9sSPbDjWdJrFr7gz0Feq
AZQ0aydGyq/f1m5wPvBsKffjIDVtVKpMltaoJp4J8Qx/opNOJG+xYInzpRWtmZSimPyZzwOFig7v
HOQ1sW4FNM/kiiXmk+Z/1QbUC13uVhCf2xLhUX1fdZQ9H6aJGiTd3lo0WU7OXiquMUmuCcmw7Xur
BXm4TCTUfqxMu8JUAMrCMxZXJyvgcnHorQwLxH+na7vMRKKbj/RtFb71Yh2VJ70Kl/Bdj3FwO1tF
f36wwdqNlnOPk2h7LV1gChE07741RhW8n/jlN+F8sY3z318p84Nswpb5pOpVGRkwVE3tUVEL5MT8
V0gUC10g6uWlhHkBezl+zJ8z9Wk9dLCv5t7TzPcswvUtZoGzOSdjOS4LNxJdFHs9iWstDGW1mKyq
eh/cV3NNOf3lglHZtR0EUDaias8vkgz2GyXWDAk4u2sgnKNPanhTQKPEw0Po5XYsr4CEGcymQDC3
q+TM9Jw9YPIUFrgIkJfShEPZapgtYWP7fngl2xK8IdC/footTR2qaZvhIQtquhJbpzWpwnyvrYtz
QOgQWpaFMfbN/w3JrR7oLBv5vTi2B3pv0i4FK1zP/5hnWX0ODq8+4wE36EUfQwSI3mLW+uN+Tao0
52R81lzHqdNHlUws3VPse2Ggvk1qgq++jw5vOFBNCQfQK0Tswye8SKZ3WmG70itAdCkqHx08ReEJ
4kiQOHhEEil5p/+U5rAGMIms2zEN+lCGH4m8ATyWc704XvVEdLhmcWXbOa1KRHh7uzbqIsUFKhux
QunbTKZOLABmQ8sBH4vOjiEEZF+OIFDtS+sVi3bgOZOLK5cbpIHb1BpNjY2d6CNuK78qkleJxR6C
UlSQPL+OpKIW7rmULJmcH8KQaU+uR8+Ie1NvkiHKj4cR7skHhTc+nhNEYI1cS4c+o20PPyyWDTVT
hlRR5+0O9pTaIGUWqk7PUWcIKmtPMdnG4LaiUPNpb7QUPf6cqgMR5SOSSpa5Tmx/mc7JoLPtcDGF
/OBGo8hjiUtH7QhL6QHkH4q/DwrsWTGrtnE8jGpDNXe3r3SjlxFDfry6JNdadVDtNkgz4SWeGFuk
MUWPOZX/nf1gJJBYpT72f1sZ+9v/loQpTJ+7/5UNnqZLCfoBc6coyzXr2xKUz05IiMcEJLlZPSm1
X6T3MMKBPyw1gJ3JSkkm9dqTFgr0p6xSD8NN6TaLzIzk961M4iEZkOvu8BQkqfm4loTSFpoZGW8y
2LoEn1SuecjahEYgEleNr2KiJoyLYKWPkqo6aCxhAEWMkluOW0oz0oDprnBGTk/7PHOB/C18KVsG
aJ1FxQqbgVUmBmQ5L6hiIjii87026QnLWErHuTPi+5by7zw69qo/LmTkdEmTI8dj6v9fVMfDSnzh
UYrNLVgGMI9QBIYHeEca9rrsqMseg7JbiWiuaK2cV7f3rl/rCBDPHBG2HeuSEU5hHem6B0MEOu2y
OIQ3LS1Tx4i4usoPUs52m6kYTW9d2Jud6rfNMNha6JLs71DaBTa3rkMqh8NhpkLQZCFv3YzgotsQ
aruz8wJoz/xcjpNZHFXzmhuB8IUqV/970/ivOJjwJecjwoAuAle6hvpijaLopJu3GhF3HSOcp+mB
9LeIijmrDNoMOeMb0jTRI5IzJ1fSL9t3kQPrrmDpFBlv73JrXYansMMRPNp+HSqyYtfc9XTxoU33
C038HwY+V8TXTTuSqATrf7QS9b3Af++zkxn78RJKBFQUm5QmZFyockd2ZlxdyyS1lGhNGaihicHu
BCLmVk1cv/OdoBqG4iAaRFq1KdVBmc7S0+mUKIgzjg2xvCIns23kbAhl8sRL9IYYMNmgRxeNMmem
PtqyYOoc9hCQesfxUXGr4tfUVA6eIUyiXylUFpr9N9htdWGuyH/CMqm1QghU4c4S0PDxOOzRcFJl
cl8kDl47BHlf3mcE988BtDcgTvdyiq4hkLlvA7VtSEtY8R2zCzQKbJT/CarINXvc/ZZIIjdoj3wD
A5q9xflSD5NFRGtFInxMsV72zJFflR7PWysQBnEvE3ng54/D+akAK+6KT4gIDYm54qVO0HA0wLgb
69UZsNmzO2Qh5KaVkUZhc9fz0c2rOhv5QVONwX9lMplmUcfzB1Oyy8XWJyszFkdDATvw4tWHah8h
/LBpZ3E8FJvqCUpz6iIgyDElmguRBMIj5Z4oDo/IMB/19GEQLAPh40dkwEx5iCtstn5OkH4yPqft
2OUZZwn7/PY+cLlhN3aP1RTqgp8M8m30DwT2eM6ap+B/1w51t155VhwgBIVhdf9bER4TIldy5yu4
pRZwwmGJfLgZe92FwubO0KLJcF7mwRL5fwrDYs6AtmFspbPPaYVsxjpsNy7nPfxzjb/HltNmbNro
fNmUNCV6vaM4075+0mL756qheLvzDyopQKvGj4r4DtLqruwdnPO/B2OSnRHP0R01dWTTtosp7bR7
xdvCAce89AHBJ4nzO7HWllLeUVjS9PgDGJB6POCQRbqYnTQCzAvwZNoYpvakgY7kjbJEVU9RZf/J
jzRqRB6PM+PJ9jhxjUL+YWdwoG+CnbLbDOmwQPl2/9kXwAvtOGgIJnfQxwRYfutTZW8YPfCem4cm
tseOR/XrNZj9wMdMMx9qEpJkwRhYojnNVh4BvDAl+/HZtgxAtvffowSZklhASKh/xynQfuM55kjY
xJyRuj8bm2ZcduUy2ntxhPirX1FmdX3GnTqzIyM+wf0399NxIfn0D4F8vKPHdjIckATqJeziRmas
X/MwMCBVYO+G2m5qRmFLPBFPaCDhjUWvYwT/qExYhAuKtjTDhAH7O0JWS7ZdUm14LA8jki1PC+vl
j7XYgS9t/B2VUi3iIew1wneR5TlfstAE52Fycgw+8nt59Z4ehG7aJmto1yqSP1D+KFBbFcTw3IgM
ucChZtkg6uzLiRZlBZD2MBaPEhPuMHQABE2YmiRnUgdG06MmQNTZ7eCNo1bykyMIMyLD2CVFU1y7
wmz8idvpJoKYMLGpqfXBa+Gf72xOq1T1O90xZil3gepPzCed5JcqOrUd92KAYE1Nr1Yn1DfGkSY1
+CrgEl+NxhgOmIzzko0LHP27yGOoDSIQTn6OvAYKcxZHrdwAFO/DNDBTAg3stoNjoBsTi+YZ//hU
RYBq/qnTbQfl7o5wrV4x3LrQm24qH10Cr1Qs7vObLXU24tMwMBlk2As0z69Heph66PEhZZK/Fyrh
mpQTvVzWBgtBgbTU9AyckggQRfSsLS4KvbAzTLfZmzA9cx23lDKd9TKDhkpc3kKOIXUJ0OzeA1u3
XtLCQpk9RLKrnaEzofOWCS4OCel5KRPSltRRouTXcx7ob3fLb+tVv182ODUygyGm+dCitpkIoA5+
UBmcsUxvkR4iDAAwkXVodlHyPGLUDHTqBOO09W1OCSSQTg7REJzAbX6igOuA3GA8HsV253D4YyIb
LSBiXsfSdbKReUy0Rd/vk8zjhNmVOBabq/ZdeFFKFMZhzt+4EVL1rHLIbcFfdyLIPVWBsiRgVC2q
18U88UMAglO4G+ha+i39pehLHdgTxZeefDjRkMK3A/jBJxW8tlQRxaVWpMpnOiwezuevRc4lr0PG
etHi0Ird6h80UzGJ+qXPeZtVg/je/z220JgqU/W6+RauzD679TnBoS/t3qsbKcOvdMlHTzyPV+20
OQRkrw1LPE9FRor6iobH6W5ugIDSHHpfIThPMDAjASALs6A3eWrey6uEXDwgfTOKLQp2E1ltPM9e
tV3hishotUKQuRYTedSF84d+Hxv7Yw1gYT3xQgaF01OvNydb366liG2JOiv8KqyclAkp/ybXjEtv
hfpGlKTr+GTtuVz4QhcjlhDFAv3M/O6QwKa8EPDYsa5tAVE1Cjytz1sTw70QcX0cR1MfFQxbyeaQ
HGS8pR9sQVpPsERanBOqQDSFAg0MzbosYmhnsU9Hc+haKG8q5gXtoGKbI7pZhB6yQfVRANB/0eOC
7FOkIb2k3b+tQm5JoSRaIRvFYhLIPbFnAbdRIMW7Angjlay9gU72ervcXDhWi7iyInLNFSnUGJbU
JSuw7dxivLJzw1YdjARyqhLNdJcZXr1ARBtxa5tw3pob6kFsDU5Yd5TVC5ZNnXuwQ3egf0uQJ9wU
90dSH/rhj5xFHgbHtBdTWKzDrE1ZpjPQ1JHsT3fvHJkzGiBkLtXmMU41YN2jHEwG/nIQ0gXHhdbw
8/d6SE1CNGCwG9yBHqgVt6TM9IZsL9bOAhQCwlmwSZdM/w9PFI17sE6zCAcLWP+9EWYmnHv24tm5
FJHOYO0HLvnJw3eSLvmiK9d/YM17lEKsktXca4L97sRu7eojV0955SWC9Mxmu+slAjmdNB5NJgh7
BaZ1rlZfgZGS+wAfv3I731bjfMBgBEhjazELCQI3OE010OeYD4M7MjUqSXdJ5ptgiIOAfW6ZAaQE
vMPr+PsHbX35TwFEgOo/nRSA1ReVos4rED1eysqhfxlY9MA278IHWyDSYIGu9QedrgHXBW2EnvGp
ze/tCVw/usJG4S/Zn3Z+Qs0JBp2B0qwNE+9eyucaDaLN/+DYilQMOysM93338UMcUrOnIxT/6upE
2q6maiqmE+4IvuntK4WhRB3X49F09Ja4TOPORXv53AZHw8cxdWqBUHAWhpw2SeM1UsgPmB7+HRm3
tXnAwkFAwoAFVoo2h+2XqtBqAZdLku6MNhoec9CDsCh9+IoW5cWTy73RJRUNhqIZoy8fFvwSvpmE
D+KR4YbF1RDHWEUDvH0HyL065w790XgmAPzlC6RI+IP0PJQ/LGZd//qLSvc5zdyHyYxosoKlixug
4iSWPutjmAXYX330T5Va8g/4dYAPswAo1SRsnFampLuU4zp7kHzZHlg8+NWp2qXHA2fCJ0srStZE
QylrWaT5w42wuVt+jrG+LZroGEADT2jMc23tbWnXeYbXM+icG6o9HpMlp/flxNPV0Igl+Hh33nLT
nrI+Fg1jW1jfq1M2biH91Qpon7+eVaTY3yny3HYAYS9sJmSf9XjM+QDi+4ZQkcN7E+tQH35U0QA/
vWx2YwbBHB1+NkiFV5FYMnIyTVnQKjWAK/1SP3XMqOZ43fHyLBMVVxshvSmmqiahgP9cWKyA6Qa1
oUF3AG/8Cp/cuauaiagwrq4tSvwZA6hLW9dgCJ8c1sW6jIEjE84HIAnkJsF0b7PDeY9XObm3/nRY
sOpbQNwjWLzd5gC/H6Ji+zCrA/JFkNBM82U1+3B936GGwiFT7DFdGoNZ0+lfP3a7WMpC2sxl1fLG
d0tbAs2zpMXSkD1hbp0RwLMCz7yudjDlzK23xlsGAPB8EMcNW7LbPGJnx922nmTPoE1gjTBEKfVZ
HsOzhu1z+CcFHIl7Byc2WG5EW6QrvJeA0ZndpMfKGw4jozOneuZEE4STnyhxedy1ZMl+Jdwu2Kg8
nndHrmfYDGDyg1weyfCH3W8C5PHVfWOVNcCDt7eMoCDGJURZt/IFyQN2ZXBTCnsXxB6NKpERNxkJ
U7U/8rphODZrFN8l+wYzzn5vV+OAh2ATHkXdbZdEhKddXK/6VbASM+vVgofLkWIMy4obvWDmBjLY
DsJiRi0TxXKql/WHFIS9375wief09tU37Beb4cSndZ6TnF81eVyZAayaQtgNwuhRbiKaMQUEl1ZV
JSY5tU5TP00+Dcsf01MKTPcYskY0Jsd4WKk63fv6ECERpaxBVadQAAV8OjQYwfhpq3K5lB4JT24n
gyMASQcWqQ0a+yEUZTD+Lgan51P7v/zRXHDTkDI8+6/Gm29Y8dQaNkDZfzVlFNidwNwHGoRFRhSe
5YQUX4pZbjtsxCykMm6mqUwBOxE1yknXYu2GNdcHNA3oa8kIl+C3dE4aa2AfsmbtRG1JsCgOAt1f
UA1y78wf2lOwppwcMosyzpDYOYK2a+hJk3oT7sSKFHEv354TNWK2wGsSwPpCoHrjfjsRyGtJTWYe
ahI7iEd08Kf9VhLjzpun0+rOyr8CUYFI4bvQFO1544Rdd1xALaNU8RCAzTjZXrS31c7QOWT/HoK7
7OhZU/IgTLy/km6NBh+CITuDfrCXQPSET7pfy0Vjx3Zippxuq0ohiEqbB9Z6gecdhd+Hyke11w/r
3iHVzQBiRrsKEExhGJbHjqlImwTfqxSeFlPmIcfEYvCD3rC7Uzs1m1g4s1+6fXQCdiKjv6iWyHh3
4DH9vZzwXhPH6IPz8bqvM1yzbHLpCW1tSULK28778l28d/TATLe3Hth+crD9Kqx95zFiVByaMclT
f8Z8VpQd6Po8jyx/Wy64Z0MTRa5lHdIwT+TYGXtozoyZEioH20yFjzh8FmPh6OtlZ4CbZSWpkHsv
aWqN1oZw4PlapEmtpsM2fzKgJZJ1cjajw0wOvL5U4rDPtU+jM2wLYCSXvXqsNtrU1tx7+CJMvayY
xzDlwBhDmhkDJa3YygyLr/vEpeA0dz02vulbdhr06T33O20cOja9vyyO5+vAfoCGdT4Xkj56Rfzq
cebtJJs+vhKxdBI3A8K38lgBJjPaB+EKFtikn+Fpz3D3MyxpfZQpEtbOsNjCeDbm9MjmNwAo8BIJ
Upv7qe33GNgVP9FhBYrKnnVPR6tu5sFCBFjUzttaZh9D7YUUUZiZI7OPBczDHRfs1BnegxGv7ZSF
VUdOKzQeNM4zn1j/Q9P9jVyWBmbJMcOoEzMluF1oypQQ03Eh3Gz88PYh20HFkTzUF7/XNpMayKr2
onurVTIT6PRCvASfNx2k6EmcD7iItnUX2E2SSAM9wsDLkaqBw6VLw525btmRG/MkzEBLO7Bibp98
aWCVv21V+tLColN7jVeAfxNs11FJUolw9F8iUkdBTlCCpaMvsYMDL+fmeQeu1c+EMzptF0yT8+Pt
2gkNxeA6W7CuswLzvkDuIv8w1kBwbRE0Wzu/NqlR88oVwswvAY5xi82pNyKEr0T9V0WlJtayyIyu
gSGccZ8Euwr6B9o9Qyf7DH+yiB0/qwg++ALGUaBfIZpbtT4liK5HB67KIV/KOjl1CAb+pat472dP
8OvJ9Dz8QfE8UTktW+SkJSlEuj+U+TVN8Wey6wN2k8nrBVyYPQH7q5B+J2O5HAy9mYAcckOfAP/k
34Ue3+83OTKAQJobpbcFld7cctyi7dJxUpSSfPRzw3D0taj9p9EmPwBuUq4DWtL2UyvpG3rEU9c6
h6uMzIqlkM4gJPE9dDFML3IOdtq97hbiUFmqgvl4zlcR8Q5yC9u/pLVeZLbMfxy5X6UUWg2bOw5B
X/WE/5dtgyTsOBdkvBY/HMI3hGuUo/gxwm8Cbjg7NgZ6JKgA9HFxc1fe1peaMezP3E7/f0ainhpP
GtaaXUruJWKBsU085ApDwAirf3oGBk3dlMkR6tQNo2wn7wpP0XF5CsdIRVzrUp/DCo+id1r5MPqs
y6ERK0RfR9hGpJcEoan4CE6Rs8YtJMGHsOZmFuIynx2kP7cqb46HR/4e8QRqNCEft1WSA3FsNfDm
48LG9xlBbMCk+4VQfwai6pSmiD5nhhmUedEGFVvAWNUAIUk/kGdQt6p1jlOWSP7QchQuXtJ3BFJG
iAP6+EfA5d4X4U638MaVZkieSVXPD6xDHOFsugW/QF1cuWB7isiDkZ6t7EmSie0YRHyo2BG50zCk
FsVsDkDYuIRvCnXwUAny8mEQ3TYrIlBOvuux/xJmWUQZw53hQ8tqFVCVI2IxfqCzE+OoHXZTkT8a
2WTgDH93fX1NaiMKDv4OiFwZx9HyU7xxuFSnOTEH0WJsrNbH+9+oDzZ6dmBAw5xanx17dQBvjLrz
qhlBicDjEKHBNQtD5Yk6BMpPFG3Mkwxo/SaoED02SaMyPyQsqFcY5x8SAG6lDhJfJygOSW/ba03f
Y+BrPI5kBFLIe+q4h6TenzD/sq/0YqzQC015EsFB/AgPOeDqC5e3fgdUax2nlIxxOCf3pMPEB+Qb
AI8IcExFY2JwkJU2DP7MYJjKiR5kFKULMmz57KucEs0dQ+rF0rx4tI+QN3tO3Fq4x5b3vXWwtYMv
dz50GHM/zG0PG8w8VbzUW/Xl3WCECJweESovKcg+o3gBbdNGXqsFhLLdL6MgJ43qKZgJTlgUIhad
44u/JzE5549T78V/2aTd5tp7etKEV81N3uL+NmJV8N22nrFdMw/cNOtbqp40Oiz7dfuRYpjUmgSW
9SbkIr8+2b/WqcPtSgK6Sso/CCT687c7rq+Um676eAvsR8Ykfzkab74lAhl9md7JuqOfdzx95bIh
18nFZ32koZTprW7kmqchxMG2GrgU4DBnNKnTgucbiaSw8tq29APF4Ys9IiTQ8OFom2r8mgNr/uz4
SuRHH9SQGnKKfg3Ojjpm2m3HcnTvB/JY4pjyoHREsL5EUw5dlhOff1lXmazJ1OwDUZu1nlV7R4jJ
523OVQ3qZcxulNosEavCRrUoze9R/1JDN0NvO/O8tjGvcQHpTL9ggBKtRVGZmd3JcdOLSIsg1YrK
O/aMC5dZdhCPqf909KQfeM8Z6/BySQOvWskPZ3Py1UkYd7M0tvzoWIdZeqehzcSbgCP80sTnbwTg
As2sERpb1ODbrqLeTdK56yKdtnxkbOAiNgUzFZH75mcL1A1MJUaGffDg/PMv08c7fiwtcX8Mjov3
/nw6wv2sU3vyycnWL8R/vgXbBPGVkxqBWPPLKlzZyQHmdKbhRCyX+CE3uafBOJq1x3O5eM6OZRB2
ZLDUXApn4qOqZj3m/uvQQm7FfSWkoYeauUKtoQXM40xwgLlhyOc2+fsQqCUeQ7vRtL6O//8vcpFA
a2DHZnQQCSy8hmx1RHKgGXcIzrf1gq3cdMb9uGorPba8MA6snIomwe2M+HAGCLaX+F+fxc6oHMOe
NfeMuQZW5CQQeWpTNyQD80ktcE8ygNA7tibtW42WiFIGSQSPnlCmpDoIQZ/ro5QkVdqwG33Pv95g
78SoM1ueJs8Tw9/Dz0YuMuV+nhDPQdejl/NPkDcp3GyO8gJNYNYmDVWbVJ2OzA0R32yDsL0NNjG5
Blw2MU8Dt2acxg/OmyVjAhs6W0pwhElZ01F50TQNACLhZ/8aLajRm10TgI1qM7xJN2AEMOHXM2cW
53EN2UbcCRhPK+bYAC24782XWCrC6Tr0d+Q6G9bemxzd5ln0Uh8TTOMgk7d2xM6pQ3rAfG1JKziX
l9N3EwHvMYADRGEbX0oRd51ZKD19Xl0ueoiKCVGoU6DhfRwROO4qzPSd8cYmfQSOy7PpdT6PUVRU
yeMTdAfGUiymhPxGMQ8QN2Lkk/6p9xBI6EPEFYx9l8rWZUAqYw4thZ2IqhK7d03pSd3kEEZdIEQv
jp2lFaYFOMMi9PI+VvC4/EUOe9Pa+JiBARRVI7Ut/zqFDWcuzdNQvuttahz6xmt9AFVQy/tQodJ0
lzQkVOaBliQrrtWjB59oBD+agvVjBFUEJo3YiUkiPsrajkot6UDjinyqVDyl8e+IaXy1LlcliTPt
ZivPySvoa40/oqr1cGPItTbSRMUnkt1rO8Mr8FbR+KqQNUKJWb3x6A7MWeiEpsjkCFX10XOmFsP2
1zYV8MmIxAKeMLxeHDZY6tEOVJusFI35jMomfuqUhXXuho1fBQ8Ju3rGb0Gup7sW6JBp9UEPoW2f
PqD4pJ5HG4wdkJuLy1LbB6j1QJTyj9K/OWNZeF3kxTlg3gnFvV1At8s6RJlN5y5GXjLyebhrHSkT
llCaXjkdHJLN6x6WKtsEARtDNcsRzzsRjFVITXY3BqkubcawmIq1UgVqcnrvt7K6xJWJuuq7cZmj
Hd7fDZ/UAkb7YeaCVj4QZo8REngIdq9aIltN7mxs4Rnek0gMApQZMm5ZX7xao/03DOx49jDOW9zx
ydOZw4KMG1r8qA4dBlw0MLugYOY90wevTLHQPjXX0DPKFcePa85m4ZmwSb4uSKnHCE1i+GX5GfQp
n2LeJ9IWYiEQ0D59ruHAYFoERKiKHkGxQEEvt5QikIXrSHUqTPjTLBFQoS7mqklHiOLMX66zInAQ
eKjU7LeuB6OTmv2t2IMLGRqB0plngWIY9UuEL+QMItHQMh5JcU6+jrnE7DZkm49IftEhGtNb0fi/
uo+Gsp7oNal1Evhjbq8phNzg8w1Kwt0diKXGGoAI3NDD0z5ZGMz/d99f8woynEReGk7eh/bsWt0T
zxLC7qzsTKnConMeXTwJrnfsgTXDbMK+cUSvFAYmRgcJm9OasuCk1Sw32yskTJJe5pUW+lY0GgJL
tU0AKWkYog5aJhDUY3nSVGphHZUA2mMCDWJGOMAo+nwWL84Xumhuxv/1V2wP6BgfHBVRqJFso4iY
qB+NC+2rdqOhznGK96ma6VfB2XdqjJO1p5UYJBQ7srXZT7YBBiNRMQ4QwDI+Qnc+n0cs1OWfnUyQ
uUCsZL2qtwkDvjAlhZUfGCClchkrgKV2QzRQu9coDs896mbiq3HLqhCJ6i5RV59KIMXXfBBl8MJI
EbFzfJNpyOjivnj0ucCDyHXtRyDV3I9FbrZJY6JgIqAYbx8MzBbrRs/TMuteHV/ompGBIdUxL7u/
CLcsWM9E7BVpGa+tQHFyt7zsx0Tlmm5k9AKkjz7P9wjDKV9blUXglZK/6jLQOcoI6mzcso4mDqmJ
aT3tGD7Mz6OxiFFhOjV4owL3/o9biYHHLqAk3ysXny9YMWunp88lFGYJ3Xwo80tA6878/qyMCIL/
/R67cR8CD6UFO6g6Cj26vAmbh1er3nowU+I5F1KmEcD9S9DmLMXEok9g9sCYf2A/xwtZ3LbcS/BP
i70DDJmWvTjh0w97K9JvNgw68302rVDN/Flv6oJrT7iQFMmJHyHwLJ2BkOagdsmggbR0yBRodwMm
kRaOy1p/H1SVIzyO6oBSJKbByx2avLycId0SEfEAtP+6zS9Kdv0gGTkO1It+xDUgh22AWeV4I0Au
HUffzaPOyVxZpbAKIv6ww6Gma4S12a2Jda+vpvoFvN5H/pWF70eB9vIAOz0aDD79RGQJDcYp+tYH
m0tbyjm+pmD9dLJCT0KvuczxQ5UZQqVhj9Gi583f+gMoIFgLESKuJABUrAzaAziJG49HXSSOAHYH
TjhYNmEAagrTZBgp7QTSl2Tzt8yySOz8u8OkE22psAltTmx6L5/wgVDUoyHzcdCGyQ75mdK0xnBy
XQWR+ZximTaF9tOLEMvAiwX75unxY8FVEE88cpJI0C69SaAe5j5NqPOvc9MlU7Z8F7HulpUfdMiT
M0tVl8G76Y5u/JB4X1+6WnOjzMArPIALGgYjhyZFzPPvEj7V7CrbY2WWz9JuJFNMUGd8w8n7Fr96
dQEvf9GwXcTSPEuZlHe4r0+uKlb5PFXg84nXVlwx43ojsnnNmtggs3YCqHZcjoyxBGZ06ni6UmZg
KrB8f2IXo+p6myfMgtUo2NjSel5Gekh8C+bDvA2M3XIwHEoeEuy2E6ZBl2motUUUjoHtmahLKmcf
cGan2g/sL5PaexGmtXx/X/bLpIPnRAKk3YwXDutBU8mP4ux7QT1M0jFK+lacdZ+LRUVrysc8dEap
rexqQb11ivqC1Q7OJI70FeFs7yG00hrWNgmJ0sIQOlx/9fNPcnFvZvHGp17vYkqVsQe38fOapkOl
yKwraE4oFqQn39HnyPQe/+rQCmBGF6Jf7EmW2ImBOtp5RmvZ0GS5pxLnH+tnu1MuDEvpkZkFUtq2
j/hzYaEVj3J88o3ggWHv+RYvsyyBYWAiuC902lLih75YXEvN3PUtcf9IMWAXKD/X87M++ZqFMVLU
C+kBjvqSFBymwcA+8z2LBqkNBj1ZK1tGSuWVKEvNwbLo58ytK2ZFPWjbw5xjVOBx3t0X+cp+BUdt
iqY3Cx3cP+U83CTl3dHYlD0qyasiCXaydjJKCMll2C7MABQ9AnC9ag+PZlVscPyWaVLYzYej1hqn
dX85ws3IE1ac2tdCltvaglUNxMAmliZ1LaRWzbmbul5cMAs+2/b3RLkLb6eA+FtfMEd3Kn7h4aMD
7spjhHjI6hsY2QFAysXq8R53htlkf9UtaNO1qlZelz7usoB6JQNpcpZH2qUeRt1prvLHMqrpYDlZ
DZTyLcvRbUjXGjBQ3GnkaPladsHfnUW+ArNIKxVkgx8OXa2KvEHuBczDCHsum8rIZ6q7P3vwPUpx
SpqDglsrIk4FunsujGG0DMZ0IrjEmFc2LYUV5gce7okQ0Pg+JIpezhimYImABeSt74l+MFiE+o1t
uH7sht/CizO7cb5NLFTiTr5rjwidVnJQ/kiMYuED+XTLgyA7Ngn4+2aNiYsze+SlrRsVoMDMn+Fn
6wCE60Rk3vzM7Xv2rmRYl7x2bE0b87OfCDExqiedLp3G6mPTxQEeK30i7eaOxPAz9j/XQV8Xfvtf
imB3GRecn4zjaWZ+KcMInOl5+toKIuEL7c3JQskw02jKRzDx/GXGuvSs/fneDLLQDOGFZTJ4N4qD
RFH1idKpQiw2NWRCdsaVu6xLVdLtAmO4PVJGA7ZaPnudsah5gTqYoJMVQ64k6/wPmoKqb6PocyfZ
x8F8s1AEf6fmPSq0jWNlmninlVJ4WhOdokvrJS3GMeIHcKgs5fHR7B7lykbq1wS/zp23v4J7IEWo
63rXHJuGyi8BzKuNoSS5hEwvWU4nlCfEQCx4BOEhbU8Fe3E7EttrUeWxwNB4Lbk2QUp1f3cNstzM
zey3pEe+kOYk5YCOVQTS0dCp6C68u8SwC7XYC9RAmc2XfH1G6dMVLZAfPhTmTOoafrpKpjsH2JFi
3mYeryC/FbtO2co7Jm5ckvLeOjs34n7z7PoyHAfo1Z6Oq5NIOINyK5/cQLkfXRpjBbMeoskswkWv
x2eM2NLWR+vdVOEnB+O9K5xNZvei0Iy+M60FW6Qzk/Dk2nho67HKl7mV2r18rvcFE0mNAs1Lw1nj
RWI3p2SqWQrYloZ/jctcYjFBbka2VaKgEk70Q2gASKUFus/j4KgbvwL11sgCkAg5kyfIV/2N34GU
pNCqyDmfshI5enPgy4VBpS8pvhO81b/PK669aG3z9aFNLaoV7z0aPNsBQ2c0TnACkbXdJ35zycdm
4WKppiAoqo7M3t0lskRdK4paj7YH5/1QSu0wxAYHTIz0fxbh/mx7mNV93DhuFGdE7u9QEvJtBk1E
aimiom3DbzAbr+bnOTQH3O7wHwpyE4mKaCt6spABSvA2H1p3YbEprKm9c2J11gVAlS5DyNjwJRkk
MENBtg2YaAkVaXdH4fSkS7/tceYbuTlag6aFV68+Vmdm7wSscyEbD84b6qNxuL0o9DJMv/+bADEc
7TKjB9O8o8PzFrNP0kO9pjfNa92bYNDSHZcEh4PaPEwRnCqRW6g4RWHJkts5XjBvsyTXNN1QbFm4
6Cowi2pKC3MpfCGPX0a9QO7Di6QiYFdZy9xLx5AJ8ELG20c/ta/w+OachoIYYf8BU9f4TE2T2PIp
VRjMe2fvktXhgcjHhEuNwhQT+vbayA1gR2LqKnHy+yJe5MGCRTOBxkBlkBnacxHVXyUNeiu3ilMs
Hm6drmvjPX0apRlBbB3mxmDu/lid8IUMhgMTAIiv84586zNhOHGISQvjhRxVSffrrO54cPflQ5Pu
hhSd7uFEF7nQB1tkwT9l2Ygfb1GAcuvehCOutfjiIiDApfDpk9QUzFvmZm9A7GyZ9+xhrG5Fwrlt
rkPcsRDyGK5GzhcrhQSC3lVEFZiQ6T7DUVHc7LRelZKaUu19XTK3Ci89XrRJog01CBAVPRr1CfBp
rdekHMZzdGYWYrojJMeUk14Xa7+OcTHBy2RB2V8XjC2T/90iMYWlDo41l1x5k2yIxcHZO2mgv4fh
5NY5Vw7i5kkjTLV5cFaThg28imXl4SvMOosQvmjx2kkvrW92eFBXkr6XKm9z+KrXi1w8pTJvudvr
uFCe+eIvVctfkiRvH6kshv37tqzH5IXDypVYdE9lLyDctBZhHMPI1GsZP54tqmQJL3Y4V2IkJ0j1
QeyF1d3D3ASIj1fsdhI3YEVPTDCO+UZroqMYATTscan2ny60FOue0vJIg5JmptahaTWe7cpHc6z4
GZqHiySrsUEuRQUTxUtBbugAtJyHhPivu8LuNKqjRYXByAyxDIUZ56Ozr1tWzl6+I/Su5TrpQvkt
DKTaOt9Dfo6hPqdkAC4rPPHMpW0miLIIxMHQreSmFqTz7HqzAUD/JZDIYu30cy8OSSIaRPc+UioW
REKJfA1/Upg4zTxd2xNT71hpvx3YbIGD9m5pDT66UuqaoTXVvzed3onIf7xX5K7OjagnwOZXVvdA
2KV3bUcFUyRstClFWX7N5aibtQ/fr2I8Sc6p68QdtSK5DUTXtm/KaswHso3GmJOGX9d0EVU3O2Qa
5wsC6EMDTQ81dIc4stwZwVV9sWGwNes45/MAKSzFyDTy03sMMb85VCrBhEol3oy+9ylwLex0nhm9
UnJ2dZwEdW4i19xHJf5uZ2Dy2vxm2unIo0JVz6W4DcajRi9mGTTFNIaG5EepCb6rCgP8cXwqMbJ8
8sDMgjwXm3UY0VDkHs6cNaJmOnsGaSeCdOiwpmT1Ct9i1cIrgALSwG9x6NHBSqDc9NyCTupLKorP
jgX1pH6ju7495AgPy7ZEphxYKL9EV1O88JegHpa5J4HNNowypQrFyvLG3lduqsTkE1av/c1fezv8
kux0Oy51gGYysxyPuuppVpwgsfP5NxfgboKmcIlAFVMT62xHmSJRBTVOaqfIEAmtPwxxTzrskY8x
zhMnOuHwcSEI5myauJJW5Z1dKgjjYfljccvKg/A2D1E+U7OZSK17CBpJUhaRcMr917ZBC9DeVs4I
gOoeZj2uV/KTki0rvajG4g3J8CpLkyuxjiMZqfIaDxuonA/VXFZrxymXFLk0yNn/VDKk3BSNES6v
IsryeX27cX6jwLgDadBJeTovXlRAker2zWdvCuj9QlWZi3t0942W3xhysiGpyniRqkiH8OOKkTeI
UVVtg5B+XD2mzGe4fDmVtNG54VdWK1Ht2iteqNd/g30/k6JUYFD2ugpRNnrGKJLOJLqn6ug8M6UU
pUJw1RzhUFYTKL9or6+Wm2qwOxAKtuMs1XMyqXH1VFrQ+vw7yft+yLuXvk4yycdCBNBmKxjpQEYA
6V8RgKUi57Lvu5MilGEp8bzNw+la0EfLmQtDOF7rp2xp/MIvTT/qxSscP1LgNAQwpopMjpl5xsO2
eQWxHWefNKbifp8hxGKIXi/Ymysfbcygl0UCgD2OEsklhq27Sh3AgIoC9PJz3GdohFveKffvWJBa
KtZ/TYv4ffCQgjeMzdHmi9MwHlV5Rz4xC8QPuPnJTTK8gO6jvyQyJ/1urZe2X9Kmht/0DKn/a22W
pO8tovnDr47lePZ8kEp9JGI5di2WLyn3WnnvGFH5ujLxN5w/h53slQ5HK1HVqGJyi1iBIaYttfoQ
g0k9J+FUU2rIc2GOdedd8QJV8Ifh9QY5ypGVCvL4WM0AgHwPJIQ5KFdrbACDTBx9beP6NQvtz3gG
l+vo5ZRe8dGPr1le1R2CHGLkUmH86o1DyfvPq79m6dexZ0iU6N06KG0nvjTxbHqhWgy9qFTRuR7y
kcac/G7KqZHGHV12NgWUev2YGgyqYM1j62kWx5ux/oSSNtg9aiNZ9mT3rhDLj8cNFPA3b9Vt3lZF
fIAOqqcYJ4wg5HtUEEIgNPcUsuOQMERniFcPZfNKzHNIOUmTU/dWModNYMkbO6MpQ9twLfi0IXUt
fU/Mk3r3L1m8EvkDEJNNn8JcSQIju8uFDafWBFFnj7VGZ1EwIa/HWcGF5Ve/iXdTGR8qrz95S5GU
6FupobUY3TQvYsd/csxSeIx4KHnznWeOeZsX2B7qZr/eXHLZwmE9yx/yDreiMRXTdbobBk1/eBzA
iwFPpNtSfgM6B5/zYIJ/FtOnWYmh8A3cEsNM/+Y0/NECxNr79Cq81eWgeOLTGE7U0olhXYSSmcG7
R1kC5tcniWZH65c/GyA3NVAU0ZD3MJ7Q4ydZ1kXLeLeTbxxOhKep5UMG1rgfCuL9WfX2OZwoJIox
lZGlZS0JFPNPuuSgDwGyGWJeRSEUa6jcV0SUueTQgE9kKzFGB0ZDcMcGgrc3u43Yd9MRGpA6YyXc
/Om1USXVymdE543L6QOUeV25ZQlTt4Ym5TJNQqzZ9EsI8UMNGYVfpMtnGrq4DqKuJcIVTZowbQG4
/h1Xm8BT77KyzmigEF3AMZpIqToL8ITXHRuOz9hO/giUqu60Pjsdw9Y7qy80+r6ELmb7RMy4BOJz
SyCsYn9xAUKerr33fC2RQaA4nixY+JZlKgZCau8D8G9NIAdC4lxixQnbTHGixVIkhwW0GN5jGq2J
g+BhaWY85rUrL9UCP/n5/7y8jnTr9OINvgTFQ3afHyOiWB+VrFRoVSWvwfB70+hz7KxFbXHCNYEN
PDMYtC7c862ku6JD6av+6BShHXq2Vh2QohwWmJS5RU9ImvvWDBT+P4qUTNSyIPyIKszC0WBLFkHd
inTOzsOxeJyeeby2fdoo2CIluqxx5IsPB81jFqEsxwadbMotZl+9SOdLpxDHVeCvoA9Id0FdR/Gq
uYRC7F9qMQIq0okEOO3Od3W9bP1HpHwWV9s+Xeo2G7963SqAePT3Klzfte8JYutcV0PtOxpm2/EP
8Vf9iTiPSlR6OlHqmB+ZqYSwHUKoafa7cPLMm+URC9BamLK1ihg1DVh3Us4wsIoqFK7DKVl0DKA1
I77kkoxWbUtyScP16UmQTwyGjX2o/tsjsx1MOiK1lpSRyOdd2pdcXO5gb0drd5zp8tsoR8YjPYay
wqRit7uklYlcqm1cncMZEpwKyYqgXOOh9fZXfsHKHWuMfuhpPzEAOj4lJ0JWtzfvIs8l00DoyTEc
Hv6nldru4iQXZY/4Wxtv87PSIreYhZiOjXgjk/RAvSJgS8wsaseqkI/AqdBsy1prPGqjEL9Sq3c7
+YcRlWBstq/FoJaSSyAEagBqE7AUWdniuMKi3I+yy1ugd3n6JZ0v+SasmAbdMM6JlCaoFqpJHx+W
2BBa7f214v221VfT2uyTVDm3P+KUmevvM2D3g/v8B6FcccbeufNDztZ35IhFYnfFYNUH3NRA/m2C
QpmYOnfSted1tbXApC4rvxbOYaQgQnxxlKCXzCq597mqkc/UTppjrKf3jG3tHd1QPoyM57JV4i4T
iaUEPgid7VTye1f7UkTEDaHocqPY/CA8LTBFzuzThESbbIGUInM10icyizZYfQM1+/gq5XeRwrf0
61MQU4YBOcf5EPBkEnub+atz+DzILLkkhl9liz83UKXmFHG/iN8Bl06cRFQXfi+uHcHcbvxpx1pB
IPEfEX1z2i3Hmijisvnf+S1aAhAskw5aRDJ+i6uCRujSY9TOe3+8OebtUlmPS9LOfyJQ9QzoAfam
EVsEzDXZc5ONakkw5i3yDZsQAcwGr8ehcKVHFqY/2VWbFpA8YUcHLMFcW1C4VbNn5rRwJUaKoTeP
Z6j2HzZ9l1q5PjKU5K3RFWAJuGElrrgnhVlBjrKTCw0p37z2Lx4m23kWzR/oMHZiB7DHcXgaKvY4
z96B1WGD2GxFqluK8WEQGhAri8b5NEbD/y0U0WoA3zL7jVAlxf2HUmmWkrnKR1tDSow+HJhhapjb
hkXtSYAZarW/YyfouG8A6je/q46VUarfMavmQhfaCE4BI6YvVAE++7N3+QdtZvv/Bhls5dSmjhZn
33q/CDJl0XL3UQPQ53+QItGO/46Wy4LxqweBueNlqu+mJDZDGEP3JL4EWsw+vyz6JfsSM8+M8gUP
z/mhbPooqAGjJlsRFsTDaLz2ITyvnjln4JiSacMvxAn1hDdM0eYQ0XdHqrUafrJXbmDGRbsfmC5x
w7CM2Emk5qQLaA5WIwXD1CmAic6Mzw2lkkP9EAIHiRp2SVxkd4dbzKH8SXmoYfOgVsHHgHg8oDf2
e8DXPlYw89Qo7ScGRWD+jUQMxL40V9hRdeGJKQfUwZbCiIiK6hAzMc91Z7chmOy2PBWrALKilfnr
rqOtHCJEta6phgVJd1oISZCcFR2ZBCWqUIqG5y2mMCtJKMCopo6qXYZnePsDk1XTx0NXvgTTWwRt
cRcG3KIT/4gTwgS0oDq2JQQhOEgyQrOupUAgo3i5m9VlxdOapkUa9abz/rY3jkSTC1ikwSpDsVi6
4cH02VcJNbVGQZYUoDymTGFihGwVSI8hFwI/kMT8muX9mfaktk+gQXYi0LWMkrYGM00bNERpkvZY
KTgH9SW/AHkc+EhvqumNI1QoS36pZ5thMU80wUz1FObJqZXhBIk5zen6+Q6yurSosmXnH+j62rps
fMbs0T13zpjFGqZf/nObuYDhS2LH3CKnB1ar8INR03G+4pPmOdNKb0hsEIFQjlmLsBHZWloa3v+f
EFSV0BA+x5P4hCzyJX6ey4OzqH6kv6s0rxLl0Y5gIKS1O/HGuI4ShbjW41Bcn+Lb8Aytx+rRbt7X
Wwke5R6ShjrF1WdEdba4nRBr2AT72plFffo4ZtEP8JNUNuv+ThwyCRA+kVvS5EQHRxBAR0AaPiT2
zhqf6WeuC86F35oijf2xil4CUjc85ixKuaNgwavgwW+5zxV4RkQ2LVyX+LTCpwCW02cHZifITFTg
yN6n0Gp6cLEfsb9mQjMyZh91EF7lEHP0xf/pS1FD9e1JADReblg7vp3CI+9f9hrSpBo4VQNPHxYM
Vu3upxHS8dSUNfuEKOzB7JiGTcxpmysVa3TSz4Oq7AGceRekGi+41IBu6gTbjsrs0jp2CRJIfotm
lqT8BpIOM2sRTVpMWjko8y9f/Qp8dwrXr9Jn16Nz3klyuZJwWQWafupNyWFBT8J+LlnQpYf2HkLI
nEq4bH8E6wxdc4e+XMh8TpFRJe4I+/un7DtM8aYGRIxCFOo5kV2cBJdSOQEho8aksPSeCMEYUKo9
1z9L17zAnxftyZYpF6Dp5l33Qai8LNEhJAcQOlDOX/1Xb7+GKJ7Zg5iri9W6P5lyuXudxXRAw/pq
G44NXa63HE1t3/XXXhsj9Vc1I2SIM7TwFSItESW1bZ5GkZCuzhnQzOju6WnC2sKWTAFV/JFE5XuT
tmekQHLOEwbuJvT/PYjTQ4m/9BRZekfwDMSvibOlcjWwFmBEaYOI1wERp52sSlegIMKx/kwe8v9s
CtRGiAgVFmeMwIUkEntABGGy6V7pYjEKFlLtvnS4aLjRo3L6ajFyj59O6VVZK3G+N0H/Wp7YHzAk
ZL1EQG2+cpw0RA1y442cmvqtAuL49s23Ko2MO20CCm9ZVX1WJ3VkKwOtqIjrurV+VoPkEreIka/P
nD87/41cba0Knld0ss32pM/hHHjs3hMOTsZusbRd/9WQ5lNcxp9ktdyZKJYoIkCYo+lKACDXfoMT
lMuuHCNq97OF6lFrrjh5BtEmflL2OKC+pCLwi+UqiO7R9yw44yE8ATs8fpCDL5gSLKXqfN0IhhZB
kAKe/KZnrgeA6ddXilgTyWxkiFg0pjlMCPufZH8I2sD22KWmWY8sNnyQFFpwS/I+wbR1BQ1zdsYq
Pgg6dZ9FNSQU8uaEKIDk7s+ryLl0LJcst/e+CnETIsrS5JJh9e4Nx701JWOJ9S64wyRsu/H2/pzJ
3IAFJjiIc7qY6WhOlWCGHWAeWWA5sKrYAKPGSjHd22M5baRjD64Ri3vjI4ZsYp2dVcCzpoIvQClL
aASjz92CNLvJUEwiwa+8IGwXrmmtyrdO/OX2o4k1lOZULTUL3Khn10MWkC7gg13MCvbMTkOTc9zx
rPPLpG8uEx4E2kR5qSaAH0pzaTjRTBJywosdci6FjVaZuLuuydJ3gReh/SI6kw+Uggc490cAbLJ1
mhSWVqJSmu2T+JTIWDtjAinxx83KYKgHmfcCE8N7UitDzNHLgRb3pHcgc413jk/zAhjLBEzpT26V
r5qN1DqQHq9uRIpdRK569CtDfXFgfa8ApdPQxSlaXsTBJuGA0JhVN1eOBanl7dWIgJB9CtH9L6NU
zwR/L4ZudnSiJImRWFyN57LaGucKaLYiD0Q33weZqrgQJzbZ2+Xpnqp/mi3wfakrKMmglDgZLtRC
WR18tLx3mF91bkr/2fX/Mc/eDNsLeFQHMc1atrFVX8IyT0aI4vSd7h6dxd8IcuLavqWrBUeHDMgf
+G/bYS+qTKGUR1mEbVebH/Ibu0JlMtJHYMeywkpXrWvHiCeMbbYoOZlC1e+piLBUuBeMvjaBVmyP
wQSINzcfhrDLCXRuwjZALoLCSJYrQz80cU/wFx0OSRj30TB2TLjzC1CDn8XgF1Gwbq+NULMVieCS
HDPq1FLpGfW0rHElX0z0O5PBhbWabhwYFPgIyWGQvyppq9dagGZjtmcrCYVNTteaXAFdbaOUeckR
JnFeqNFczhGWTIlMPtr+jCtJIUloLvCXhvc3G8B/PSNqEQ6PldaJJefwdnljwtBLKefvAFjJUvGM
L3okIVrSJhsnll8xWwDtxkSZbKHtqInzUBN1XMjqSSWZNCj3u9WLA2S6ykXDpo2n/1n+R/S3ema7
otQVx6QPWXybIa9zrgHub7kF4ahpZLTnpE3yacVClPpAVG64ArK6kXiOAwH4FgIiZ/cLzWoBlR9S
ClVxQA5o0gJzDdUPKoCbFPSHTMQMirbFXA092Lblx1G1Wzt2/kBAaIMIzIMhFFkHgx9/STbTCSev
qPdxC8b1dL6jyOGePPwbbmAokeHWE+APrtHZqV415J16365/EcM2lq3gs9TycXCqSa41UXvqlMnw
r92ZC/QIiuf8WURnl7uKAIjJ/nRuaVNB7+81uCnRiyOx2pvGeoh44FIrFG9GY+ZAK8xtMhoXa0uG
Ix1ovyZwj3S0mqd75KtIBAP34m/DW7q59NihsWjbsEKHZKOSD4OHJXScnQJDZUs9sjNzoDVbUCqT
8AR/n0RhkdCwSrCem2PhzF2KRUYDMK+AXkSKMbwbXrLqjutLz+p3SgSUqSD3+2VNeTsNMGwQ4aQ2
odMw1nVNr54bYhnLccWw66naSKLMBASfYtJdbmwTKHY/rlRonipUwpG1Lr2QYW6la+o6hG+dFLGL
OkNW0rB56e+FqoJgNLIHsiIf/FTDkFk48cd0/PJQsEQCHCUt2IB5XeeNUPaSGkbXUwV6iktdHHu7
L/DQ0iO1V1fjLRsI4XZvj06dQ7A6b5ZfvlrBKb9h6Tz7hIFcfMc2Ndx6l0xmxS/keHp2yTnJqPnH
g67gXkP/1EGD4ptpA/NUL/gLIlMQhe4GaNTRIRFp6AkGdWJkRV3SHXlIw++4jGC1+iGi3TJgTxLC
p2/bsuPBhjAMIE73m7+Jnt/B1m4BsBP7oRhn2sRE4zhXCW3QA7I0NFCbrh340a/SCZZ8raHrXIuj
8DKxi7jPsWJHh0xQ+2tux/kGbKsiAgnuywaugQ4187DJc4U5Tp5GUliGmPuxyOl1Iof0ll/2uE9b
Eyik2r6FGXnXvxA1HD7ZGt/JDMh2Nmj1Vi/IxOmfGH3tlC868ZzEaOKVC5sRS4ZAVz8CshuLhHpN
fB0P65w3IstVsdHlx9+MKtvuV8Th6cq9cODAyWu1ag6xh3ByxUBPeuq8rKEms2cwikidy1+220dl
iHNEdbB9n7ExKiZwvg6ndQPg1PashQeDV4cbuqIiUOTb6UfVffe0+qnVLvRwogG24fciI6Oxs1K9
cz+hiFCxFAt2BpyOavaHvGWrXTwHhLEKuXpCMqLMYyn1noaURcnzvcce4WuNwDebZkpZy1JJxMCO
1+M7p1rdle5bpwN0pkpmvZHqYl403zggnp0m34LPtnllFGnbFMUMngmHj9G1mbnr1NAUhcxR3Bnp
a4OJToHKGd/EP/dGh2RJ9uRSUG4oQQehP4HmDm342GZ8vipo7OIyXJgHVJgnvDV720643I3d1IZH
+Zd77x4gnF+M9fUHzqF2PQkJ9Uaep133Ie+OvfZlfrZ9iXZZfJFehzss2ApO7T36G8+uHtVuP0cY
zEBJ8EIPhC+ytDjnTI0gM2k7prkdXaDjowkJr0/u+RVCWB4SUJ2bd6P2NZcU0dx112pkkSX/wHhm
L6wwgAGehiSCB1eUUtiUl25/nwKWccbgEYrsUUtZeVTe5A5C5wSU4Ys990oqktXrxmgrs+kVlhc1
GJ4zIF1wtabCV4BALjhN8OnefsIiN8rLmSsjgT2ff73oXrIRb474S641PtAkBvz4Acd/yt6EbuFh
GcNX5r8jv4MQJs/cZ8wBrFuuWxLj1GN/QMQdRQD5rt65tmIuW7OU+eAtmey3DnaIWmRJe+rP9hht
WYZJ8iHHMsx4IwPwvgyMGihESiLnVUOmC3fdTCflzco09VnQ+SMUWIuGvVNgOCuVV2jT3cMGg7Er
N0Acj4gejD/cdH5itZvEyxDiJNTuzlmMy4PwHj7AAas1GdIjbITJUFzgbKUZ9wgbAsK55LXjn4/x
DJoIKd2aWlABvjbz2WbVgomOBBsZgcFiD35aRj/t4jwlqcf7IaGmI6BN0V+DiNGRsgTLGsC9eltB
lPoYHQkuvq8MfjvUfIMoaBVtcOLsgVAW631aJrA1nUOMuA9lqVJfk110nw3DDoVa5f1l9SPDv0vn
evYRCh9Fi67noS8qaEAg0BaO3Vk9fEXisquk2y0yOjaaTErwsAQ+YR1q79gJ/bI6f4U0c+DVqdjW
ER9Xny2YZ4UOYnw7MLmphUJfzkXzf3NTMiGeecISHfYfqWbFkK7TKa2HFSp0Q1HyhgiNbuwn8sGw
kcJalkJxwrrqlzDgSC09VVAgGy7ghxD4SJniXpFa37YVZZkN1G9oZdJc3RDwoo3t6707DaWaTZI7
otnrQSeCH0Upq1uaYqMaSppp1nxr+tqY8gkZAAsdgeTB42UOobWHVk/q0i2XlECT38T0Wf+8hoB9
3vvYsvLdBzmMNG7HLiirfXZQtZI8CKoUwM8BXTzQTb9BPacsAmxVNxQJAgbjNx7WKvj1cBZ/i1d2
7+DsOfx4cQrtinMJsx9pmtUMAIrWrfuI4JUf73wOdF7coqBgUMo0UgL+kN+Wp+NW+FEidsEs7Ge8
AVlMPUBZvabo9di6uffh53Fnwjd8OHqWs+4WYz3Js4PXILjN0hxA/idg9PPnxvRF1c73L/3ev0Tr
b1IdGnoWqNdQyKZ0k8kQfu/VFaHkKuGfGp/n996t8xxj3sNE+SaVd+9/hfIkDE6n+gz7UrwHSVpP
LHqVCSp45UcZvMOUs97y7ZW7svupKHDDOmQWKHn0/0WGpPRSoQr3D5Lrsd9kOHxetDm5JVtN9cQC
BLrYgGat8QqILn0DHPSqfDbRO6iDdLqvXwBJjg1t0SG/wX4ErzY2Ru8K+Tj3HQZ8bL4PG5JyaYHL
NXgtNlOFO46so0SnHvyBzJGbZYd98Z5QrdwzGSxvlmNVMa/bN3IlKyvzwdN45c7rHGvE5zQa7F4y
U/3lmSkUPkN8hCXyzwarFO16Q2puKmr5mOLbUP9Bnpez2nbfkH/utF7kJafPBBXTrb3lOwuTZpWi
eu1OM5TVzqD9H+N9cHDoaHD9UODyzpGldYIwlcJE+A993JWZsVYqc0vP6sg8kkqXiIqIYTiY3lNr
uwNsEpZAt205Hho+ogSHMGmRpw+IPpbomFJ1rdkBweWUVgbfm8NJcjx2bTOiR4kK0I4hN+7mcz1Y
14hVLSlVzhm5q1iZwvhRvFAGnVh1zq/WBqBaf+bXnbd6f9uprB2o38IOx3KpTtyL9tIF2fvN0MdX
wr2un+H+sVOlvoNNItmn+gRov4utpWEjHVSLiQTwgG7z1SprXqnPkRxKAt2Ta68AOLIf7OIXIiSl
Ru8LQeEvskIkMAcu7T/+lFejs1dYglZqYDRwO/22b5ea2tMySUnyMO6TuFk/cWd+yBI7Ja6IMssr
cMpZMvaGBI186bQmc3PIP5CDKy7wgf5HbhFOfdyJ6fAjCnaCyYAYqw6laBolOFlmagvJX74Lw/qi
FEaV8ypHuPfb22Qaagiw9R7Z7sC2g+uYBJY3aVt0yAvizQIV+fYoKUvVQZ4sePtbK+53qKFCB3e1
G7JGdiY0OZZLl60Mo0oMYb92w+JjavoEHRwAWY4/wCktsaj0aVEC7avPG7jsF1FO7lnZB+Oo1U2/
1Lt4D+TdW2pOO/jyaDgbDP3ijNnLQ0zJPlaNvLXsL/VMIu+Ne/Tw9K9WioxlvjRPR6fMQyny4Sd4
Nq6latOXuW0vIDTuTpQFaibb1D0i3PGG5xg/D3QqvmauB+2VVsrarSKqNlT9TxLr8wMkN6XrJRra
cYgb3kWpn8FgoYMhY15EGTZRKCUTEKo1yOe1Q04Hzui3GMoobyi3OHHn7MXXqz/+s3q+yKoI+/0C
r7HjSXPu1EHXNJFaKfP8NgQn+ujfDvvoHbPUBnwYwM4JQ2Bfqg6796acTsCwHBKi2OPDN6zNv3Ny
8Hzj/PyyTaAd9zDKuXg7cge0lJn3PCkED1k1PC+s9/fdl9x3U9NaZzS5GjdIAvmhf5zDlgjLvKIB
Kx8sSYzhz4AUa+lgfuz9AMeNRcS2J4MbbqAoXS4UNp68w8tpiHwf3iTMtWE3ba+Js5OcKGf9FJYC
MFYmlabXb3niiI7cWqOjQP4KNIalnvV+XurluU87LkqSnLjgKcSM3KqEvH/39MGSuCdeUSNqh/fH
/Ut2EyuLs+79XuNzp0hYZPpvZFQlpFDwtr0dMM5pHn9L9PTTfeTPaSsJAR5yBwIiEFVrTnTDV8pX
+GsovRjcG+tnYhwt07SJmeNwaQfTHnNiFc4rwnxhk8vKnRc8CkNjZMgOtvfBwUv22iAv+dzBYlF4
psi/xiE58mPigV4vgynont6OLfk4zKpRUamMwWWZ2ISnDtnAQSpjiz7ify4mJoqlU4mJ5eVZJcFY
kBE/Aa6DVkZ+ngMccgMWrqao70ziSDQ4onvNfj/qt9uO0ge5cx+x2H6Tki/NO5UYoDA+G2OWmrXb
0vEcLFa+yzURca+XMH+45B7av2JadlqBsw1UOvy051tHz6hoCExXcCAIg57frF37kjp118kRGvpg
SVH7pqNKJSHuO7pZe9DrC6puoTAGj/Op3iklOtn4n1YC261pcrUPaooYM6xncMnam3BXAmFVLQaX
dh2SZ/jb6RL2hVhW5X5oH1KCaILbKFGA8M5y40so8cgZK1RvL9ol4dO0noKh4gjvr/JYGzxayOIb
5mBx64kxokG9NBFcirT3ZRZNyBcQNUv6GgFxqe/yEOouPWjYfP/wdvmBtfkReKShy6CkVG/8o0/u
3lWmnurHV0859hHDllmASqpUyr88oiYaSedz0hOi9qekMmtRBAnSgevjs2NGlqxgwCR3NKiiyoZo
tUbuO6E6P8rcU9Fsni5idiD3PlfvZ3c3RBrX9ajcjLCYkUswjxjrgc7KhErCtothCuCywYgA/5xS
pn7MQPQSBZNhBHWyxsksq0G84zVdykSIjoRDLnp+pYH5hj/t/pJMPhEMXu/mI+pXRh9OQI2mkD3q
QaYpSszh1w68ZmgtrUstgIhDWoDedEJ4aVXKermBZ1UUrSSQiFEyj/OnWyPKu1IfT0LVO0n8zTyI
YOz+jH32pVoXrEIwSCsWH5OYtlQEZ75zPHEGfo1wUqcURPEy8xjMqx7gTG6Qic8zXQUcGl5Het0U
AeyOxiUqQduBvUSs9p0WkzHXY8mpFteBkg1uD1giLIb6HBW5LnVt4fKccLfdtBqqPUJ0w79rlmIl
gG7yRJ74oE9QAyIzdjBl7DTJHRU5GvmFxgasTprSE5vGS+5jJ8jbdw6fBmwdLn8yi0u6KFAY4vPo
C1jfDeJHz7MO9kpakDuY52WFLiJWr6RmwEK+cWLclXSQeGs5Xb9gamZzvxfMS5c2+ndz33E8SsCZ
8bhszk2AZjQNErJsYOZIE/bPBKT2zalpsSX9vzqijDURVYO0vI/rN1m/kVp5jXztI3f54D2CikCL
KJF32BFYCYfOtLxoN/M2btZ3Zy7QlwO/MfjQQiEg/JedVQdCOxfEncHm0ohuJstL9ueAgFzgLv0R
CyNd1sf4K8RvgLtpOIeCZeeeTP3z7cRYLOMKad/pb//sq649UNh6ZdcprSU5BzcosxBqf3EeJQqC
A3tweOtSYg6rWKw6crMRN6KOvqQdZNsZQ0BltnnhAp4pP3hp6XH4I5r22GGR3grsONmA+87wDYI7
dUP/5X7xKqsomwJXdh1Ah63sjCWeyYD2WPJmEuNTa/vw3AnHPax2GFsqydTR76YNHVFJrZirk+IC
4WBHZ4m6QV42NpFHtXyajwr+jqnXSwLrwTk2SzFnwcWKNEtgvoEAdjOz+rGkWajrdadicPo8er/7
FLKTzqz3ias5KrYwdDYdHfFPJpt8Ebos+XrJiMRK3xvflR/CKSBlV5kiJAENooOeSFmE6PD95G3/
aXV8VeBY3aYGUy+JfUq+P03gLzbnktSzpHps1Rhs6dcGGlQnoRbJhqMJ220yankQ7x3iJ2Wf1wi6
zDAfZDXSEU4OtefCmxOiOmLGkn5m4r+juKRf3vtJhXnzSBCO96XUPkNMYyeaovTvc9TmFrR5Y0nS
3JCzw44RcE3prp9T5CokAkK9/a0cEfYXFL8sQGYYmROrNxcoA5D3ig5SljsHMkIeTvTNZ78rXzLO
1qT78mKuq9zOZ3yyvItpSKk+NUzr8nsLtzghayJ3OgbZNM2ehpyPT92A3RfMOL4u5R3X2CydAElE
7tGpg3ttHNkQaX67HuY8sSIqqqqABA1iz2xYWlYsnJ/Yv87Qzt2UHHTlWXiGkxJJZhKz9iJDXPEv
PjUj9Y/dMc2NqrL9JsDPT6Y2aGzNjlm9FxEzMBpRmIaZNfTHMvcI7VWxp6nroxzEAlmq8EtR4NE8
6rfAbgtB5rlwtVFPPWh+iaO3HtFM4NLYCL2Ge7meBLxXxa+92yr4Oz+sj/GoqxsEP6I0ZjPD9MO/
MjqPBhjwkReg0WKJ6peCZgRa+DsIuTLqo9AnBS+ISXmeJwPyU9hSlM4f2mpuLSqFXOPaGYgIVR7N
A59vBUhWbTBfyKAC1pD/ZGa16pwwxw8erN6i3zn0buzgTdvcSLcLjfPBZibSk1/MmkD/maVIy9K7
uJtTe6dKptqcH2GrfxzyQ/gVL+zP6n3lbYu+yuQ5GxpeIuwFNcbObtfGwjXNOxeCTiUrQL3rPTnB
uNZPM0DunDvOSzK4vTynzI8Q2c9cEuJxP1h5LAnJf8pjmZf8r0bsM+LGq5rNNnKqQWr1oCsjvF2I
mkm5TVxT29ihQGCpHwRNDrzr2cenPyHqJOj7hit3uqUc59J5s4zMkKGHdbf+C+MbQeXqvl0Dc8Ke
sWvSFLPR1TL70/fB/Y05YXDJkBxau6Qd2glshFgaJKimHH3JKlWtsH26kth9dkrXk3+nrsWrwp/1
EgQujhquez2ls1wHTAfGyG0FIVfDtp6CeLENzYRVyruJi3roXDe25X3Xw1pHW129ejPxvlgFu4Mq
FZ21ONbqJ3xN9nHYyApXPQCM4QtDDUzFQjbz2N6ZrCb6PA7KhPeInZKCVeqayKpNdCwmv0UTG6jt
trE3Dy1o7Gs7KsVCCC+0WS6l0gl4Cze/K0JuCtpfwrhUUjdJaA/1m9ML1pf7XCmIpr+OSFCrMqIG
LcQkWo5pmOxMbepc7++Oq2p4aTrjxHuZN0iAAs1x0otbCxTkmtP6nRvmLgUhAwmoZXL1hI9/+sK+
rAJ9jnHncImnPYqwvrTOs8P2CP2nd7j0RI3Y2PH1GQZUN6KNKC29O/sZfTNsgB40kVMrnitE2/lm
mnkZ2g2ch7jGFmWUQIMtPDSrgqeJNgoPpMWD6Zqe997qxyZOC+gX+Pe+zbv/iUduVpWmP+YkfHCV
Hj6XTYBdXpqNH2mjs2SHhhBRgj5PP4XEosELGtZclBE6viHddCwA2DiOiztceRU5jOF2qMspJY7l
vHYpZW3AT6QHfh/uHElSoYAsw+q1+2LllqkpRO4a8h1jc/GeiWGNL5pt/2ZI9zwprq9tLIYYElg7
9EwYil8V+OsAMYeTee3TbdM1uihRLZXn/0wNVwIlrB7YKRXzsLk/E0p35PTwVvRzhcdtRGXeZ/IV
VEsyKmY+X7credNBr1lw6HG7PHMMCaD5jD5bXdXG0nFHvCfqNYskui0a/JIHEl0oY/vI8huQnEwF
wIp7D6xOkAZneRdcHaxXDvPRNZAT+Yapss4MLBOORJUtYp2GCI6PuTW5jwpvHwWHb8btgGxwiwOb
I/umF5ixRTHg6sWNnEV5Gwv1Zwhpp3Oae134IQbPXaRhlXjyi+afA6Ab2gcVssIOdGWJkrT3jzaC
IXiqrYpgHsj4+Pj+nwJsfyOvQRkTmEh7LzKxRCZyCs7eSvBmpUSsHwQJ3YiNWUb+qk23Y+FHa1Uw
RxuzmkSAwVWAm3zJtc1dHbxT3XzXNt5hx0H+byMq+V87Spx4oWekkWnabxh0E3PPnnGvXhEZVMMR
bNOKfAYR/glKIBiKe+F6B5vyIX2J8gbs12KFREQ6JlGk4MjAp/gJuFhacWSF2/nwLo9TPy6cFeYc
hyzmKnjR/sid56dYPp1Ajd0AwzArxN3fFUfdN11uhaFrrXreZAWJqhFBpMnnlXDFba41XMYdHsk6
V+No+vC1/kuyJZwk2Vbaf0+pBv/RyegmYyZHLyRKKn+rV9NLLw3KZMdvukDYJ2ONpS+gBx5F9xtc
o6DqQA8wq00UyGTk84nm7iqgC9vkRGjwvjMIwYeaR/BsqlaKajgDGt2L7GqgIFZxObJPxcqd8kVh
KLRl9n3SNagYsvxjgBX7rq7UIw8gDJRRbrK6vEYO4/7lUmNmYoe55tdvDgTDpMslMxMACsueGdN0
GAV+5dbAypoT3JCT9a9vgApHNK84BymlR0GwjKvH4JLaXbnOPxElzFU06bHXmMpCoCMKQeiZAMva
V6b/n1f38h4UElj/M1RKSH7U+INqiAgobvEsKNOTrWDFxqkpk/Ov2k8mAh02CPQRuvd4pmazqv5k
puYHfc/suaWwNddFKt4Y+FLN1+LzlepH4sMRQn2LeAGOWXnqNZQ2bZ/U4WJMMtZjK4AJqCxdk8b0
4vKq4YfaWawuJLufp9iFBJuCVXgy9dg7MRITvCHIGMOmoBEnwDS1QMluV8R7DuTA6w33kOKmMCZK
8YODjRz2qvcCFmUf00xKqdd/FVY+01DoVIZgEpq/svae11X2GGQXFbOFfghOmZstuwxtUb+G9fUT
Hh2h9c7zJcOkZPycToFSVRC/iTAUpy/TBb4fnEPnVi7/N7SO3PbNN2tMKmWoDkaOjNoRxC27vQ5a
nQ8wqwbXwYVNjgjs2axiau0sVPxfyRDiMcGS2lIM0rLneX/FrYgvDwvTVq2cs4bFwPh7IQo044jJ
UR6apcfhFdFq9mr/y16RBBVJaK9646nKXl6S4+enxPsq2EOCFNlpW/snbLoQhUyhrbDkZ1r7QPdt
HxZPPH6v2eWStZi0MFVceicAvYJywUNIh9/myqqVAyLU75GvMZMHZAFduZfiW2L9QYdP6uL+AQ7k
9JvEGf5tPrClTqMbw6hTINdanX1WdHaoudNzcOqZRYHmklrhqgO0XfqVEwg54k9mLPIhH4zwBzWU
wcCfIZR7Y55qKGfKgjQTLlLqwoDaH3bLpII4wew7A4YVlhy9S+H8xAIZcSdrMfISttdS0ZQLrGyh
OUH7N8MZplOyrBnHSCK4mfQK/bhwKqYSQAtCmP7fRhmmiV6kvx/hjIyhsQ80HpnA7zFZ6ndvawTO
ot+WI4MK8n26RAT4khrgV1oEAhNrsXDwf4xqi+kaXgwkTSTJcwgnUcwWLGizXXZ2omeuBFguiR1j
M/JnzdmI8LvrNeuJPtNHKXBJEbCHpxwtlGtrkjUuU40MHOdAbYvxYgPECvIOEj2s7FzN5fxbNAAd
tz+kkAlqED6l/DM/ZQbuLk/oSx1dqPxr3YKmnRma24z6zsU0EkkD79v8v+pDM5ohqOuojCRJjWMY
cddcoJ8PWKeODvO54+qy8nsUzkBPpDsJjCjo3HzcHecMJnb/Xwv2jtkPOEOL7DNVVlHP0rubxp8o
Bj3HA2sPLnOIuDlI541nHYVm++iJYBVXaik8pdHEv0McOATy7GhdE2weDlS+oHaBVktdVDc0knsg
TShDMRPAzkeeuwJQXGnx+kNlS+SS/QWrPG92Bb8CF7fSODuIwFqtrjWCId8TVXSiK5cv35oScnAl
q6oqya4iAbYhf8jGld1pe3Ee6EZHBdmgCPXakAXNDGJyvbOi4qd+scVlocLVhpeJZ57JzEknSF39
XAU/muUEyGDZA3vSBS6rwtm2eLXKI3bjQr4twdo9z4msvObaUso8gvzV319HpLRa6AE2krWAwc/2
bZV8fxv9X8wcxydwc9c8XKnDX/9Wl4zRAFI3SNFwHaw3/6L1di/x2dsefIQbH9rv1fFOkNY+K4LZ
qvf8Q0PBo3HaQhhFQ/dBER1TdqvKsET6nEmb78B1yyI+0fmHSv7hixP/bmibHzXDWLqvvKaEkSUf
8sO5k4rx6kUtTOQMv2snBI9avRg1LulXjHqPqCK9G3K65RWrRO4baTzdRBSGJXexQcmenriWsgqs
NdG7meCrI2GsZcH0QPOd8UxiXAUGumPZS0/emb1ezaVIQgQ84SJoLkU2FQKsKnzIo2GoK3YQ2lOv
/OqFJOfmYKIZIo1X00EJpYfBHkAloQpt8c7GkyMX9J7YqCY3tQAPE6224/VypxglsoYqighh99es
ytrRJAnIbc7Yg70efHLu704qRY7X54ULhBuf4U5AlId7FWg2B05SUY9GNNfGyblFicjIw3skXphe
7Sba58XcKxyLLD8GInVo6OgABsQwqLx89HHMD63wwE7LpY7HBXD9PiOf1WpTbjMLoZilqHZ2vY+b
ZwSxNIL0RTMLcP9o23fWVwagAgVylaTTMKtcfy6hpExuKGPWcTgIYgUuo8KbXjJl3fJoF5ex/tX+
5cDsUbmAzgJqYpq6hGsIb5QQdOiysWYfhRdXl/FV0VhHom4/ncgFdORZcs+5ywnxmVOpJwuCo/AS
mPEyxGQu5PThVSwIZ0MfAyJiwE733EFegSbblcRMFc0c8RfczV8mzmnt+ML1K+4sJ7EZg3riE32Y
1Lssk43GaT5lJL/ctUK9JD3DZgcTWW9Q60qHgE6IoTcoSHT/W+7usHG6tb+mxwVjGTjc6Ubq6kV9
qrRbtGwgetVw3Kicsfh7kmRPLdbqcuC0zNuv3iazP9A2Fm6IMpr88LsGDclInGOpd3c0LzMVileG
wixgoWmTVK7hpywJB/9b4nXBed2FN9l6r4mEfB13e+q+bDMUUxdklvebSIuFC2yG+IGxhcA97YeI
ehcrRs7Ji50XI6yhboFr0DLhnixJlyOtCA70W0bCVXnStutL+NVVr/QcfD24k16d2JoaYpf/zg49
HFeSzgdgvnj8VG42adPbRLMuWbKHV7o3btuOFZ3sOigu53f+UtQNjnLSkVOjKjtvelQgu7c8ESWT
s6M9hH/olodSmCtsnAGVB7h06ji79ru++3KEqf5TZRavBA6e3bw2NCSa6EmMFa8VdJ1xkmb/bwUV
JdJLS1sd5Qjhb553luMhGZVyRx32ONLsFbqnncM3BVT/eAgfhMw319o8SHd3x/ikVCQ49KM4xYA+
cVrYU/9H4HNPmC+I5A3iyYAroiFZ5DJw3nQ1RhZ4iXmJ8M37NKibQ6ATQGx8upze9z6GSkSzDAE6
nayMjBZQr3N9lzbOpAHTUrljS4+cNTBZnvST05dtY9J+KM3DfEPwl7j8B/5kr9lLi5Y333sMVBbm
fxygIdcUncnmDrOMkV7D/E7B5pT9PnhkIEQ2JOcC3ibYkecc31KUPlqELN6F6DJkHi0Lomx/7Qrg
+khsB9miWfu4V4ZjwJx4JNy+CC474OaRWEFypIpiA0erhtq+pCzOQDqV/Nht3wA0wUuNvLryl1/v
/P+WY8bupPdQME7eYlbi6iDOS9z61A5IFOqYMl1REK6AREQbcILilfMJGzVndmBWMWa8zC/MCLQJ
OYsRISRFx/1grf2r4He5ISxnMiSlK6iKK0xQ/Qcu31nQjp517dAlfLy+hU3j+kog2FXyGB3YDMjr
Q70MS7m9QNOpTZ8SsshMFutUIugUpvSal0hSsuIJC3YPBNKQqE7zkyW/sdgxe5mAmoIgD+MGD88n
Dr4TNVvyVoqKELFx6M3RY5u83b9Cs6CwQ1oe7Oss0MMr0zvLZEm0NN02RcSsIERPaL4ZgEa2XF5y
fVYd5/v6fhBEm5lZq9tDeo8unumd+2+0+VtWB/iZEAgQb7oZaQDk9QB7zt0SjkbBtd297taDSJBf
EFqwd6q3nJyW7R7i51dt2uK0ePntzjC7QamTqeGEPnvoK1Rxt9uQ3Ez+xJ0LsN6qLpEv+K9NTKtc
p7n6ZVe4PiknNMkRPQqSFAPZCsTmPsDg8xw3gRDiyLKVQzO/s2GolK8pk2sn/NsDsfczIzGnZvKX
1kVzFtIQP5W7cgInVvJgerYsV/KSIbJxUSzOW/Y+CyNy7hyHUX1SOdqz931Uyl0KveFK8j+guvAx
zz6hjiPmt8LkjJRVxep7K4YnvdRqSm6P4I3qKMOC3jiyoU7EypYZ5QVZHFPCddsLsH5NHuxpGH3Y
T3Ef2sFEVN1XNI2g8I3ouvEEHxSKD0/7NJwWekZ1hdNQvWXCzrQoQ3PqoNbx1vw16xR4mKQ9pO+I
dciV9NUbvkM8ssN8IoBg3F7H8j3nHRetBxVObsSY0TE7DaaTOQMDkzW5sOiK+XYHsW9unZfCaWO8
nTFxe1mqddRrK2C3t3cc1vYxW36Ih6ZDmd2JrQ4tfLaTa2tZ9xx+Pe+O+nsM8L0W7yBEIhC3+D99
kFYgLrBIbYBsYSlvNpvKsN8rtZxBFd0D63ilhAIQgBYf35QfGr9fj47NQawsIAbK6TPaecK2nG0X
2uodcNR8xT8zNGRcIi9IhhgvAIRh5XFYw0PmR/CFRhyQHrUw076MBP74kzVr26j+Pb3MqGgMe8uo
RVK3ktDh05TxJSH7Sq67Fx2xyTA20suLjIjeDSlpM4IXoAEha5yq+O+urwtxVBY7r/SlmoC9THZ8
VKnTu98ekORWuU84za9S84p2FgOlJmpoLIHtenqsiVPNyrzJ5aaw2nRzoEn/lhVc363w3D0w/WY/
IQeUDXxQZv6oMudvO5bk9i+yUahXtQfnCHEz52Ir5a6ojWXBlOOW1Nklu8I+T+5U/y6KD4jtaqj+
xFYJPdaZ4OYEjtAvy1Jwdz46sl5XBf64KuJBT5S7WwQO0hcUUrFZNraSkuzpjgiA8aWypJ9qsaRr
ztKfaIYfxw1zVC5UHAsBe1+AfOSjSWD5nr7Fun3qFUxCIoqj/6L0nN7Lr0hoMJY+MjAtJBiKYiUA
94u0NYqXduK8h6hu0f9AtQZ7iHd25ekeFy2C7CBOys7U6R5KylinyRf7dLNWhTpZILCbj9jgdVey
y3Ye3Z0nrrU8S9VHWqme4HEsjLgbR2nDW1s8rMhHM09sSXchEoVbV2zZXbl5CqdcnUIGTneRiws8
abhygy7l2131nZh4u2lQWHAdTyFVwwJ+IAGdkROF2+tSL3yjNixaqncOU6FUqyoF/s4rsoprKKz8
jprGWLZzytlBwD1HU5NEXwRBLssVihkr5SubPih9PpNTgmlRSVKcmCGfJ+A3px6IaRajtx3ayot+
CC+CZGa5TVmCdcYco46NiLSjKlJly7ZXilpVTxeO74iUr/WH9eKUOIZfsX+acF4X23cey+ke4hHn
og3oYj7BxKhu0/7/1AXHUmiUIvVjVEHDnVNxXtct+UNJM+03PGf6eDwgEF8hFPJedu3S1tdsEnah
wWAwMym85jLUbAHXV/Gbh7kxLP6c16q4cXOOv2SCcLSTP1vpp3jRC4Suee02YGzSe3EcQrmOvq8o
gXzk7YqaT7jl4UMp4qhUjUGSQlXTwfgO25Dfk4RULYuVqSH1iBjpfg8UAYLs3OO8y772y2PArcRU
5k48UbWk7Qu3rEqDuo4PZv+k3f3OJTZghmL2WkDEzibK/E7lCZfM9NIqtQrdY+vQgc3khw5tUStK
85ma/15q1fiBGcsHxW8aW+xVCVqqsAtgMe93xPqw+p64YH+fI4aqiDscRO3RlkGTH6ND68wPCX7M
cSLkwzUFhaY5oG3XTXNSJrBcXRbvYvpHeXYNVm5GR2F1LVYShPJKirVs9eCWW1p3ZXClksOSkQUg
VPjbx5zXQK+KFV0qAjHXPWpEhGDIY8xb8DQ93HezV7l3AY8YGiw6C4FJcl85fWrduPxhRuEd5x96
7fPGv3Z+L917WCz0CYS7fDgRrT2mQ69sdfpOiDC3ZwnFu5TPBGkgv1sUOs4ZkVCtD2l2LzhLSZm3
8Nw83Z2UFXoUVnG4ACGGCgPJozeH5J2W+G/YN9IkCKlzxXKhHjFe+V7JG0ldDiBtGQ3xdyWL0bLn
xKlylnxncLXgITRR4ECtMjBcBqNTIrkZv5rffJEBklIOPf4mzhQsUnNZE/kPHIIFlaYtOMFo6pD9
IN6eRfoZ3KuuQzIufdiA8V/82Yt14Vg78O+fY8BxObytKM8wt15Aq+zxNbeonnbfwW1O2lZ/7Ik9
h64atc/0wluRcc9qqEqOc0f97M9Ij2A0wpAZkKrMoWcR+yD3RV51CIHkAgpghZVnQ6m3d/OFIBo7
/t2NAw/Mnw6pB+HVxOPQ7aQb3TQxKEIa2HB7GHm9/VS8gNQCDd1rxZWPRN0C2SakMBwRsrNF4PJZ
UjmWGi19l4vdOpC2eD7k89i6hl4hcoD1jwl6uh+d1JZV4n3fQVUmpO/c/MD7GQuw9QM4R5aE9IXF
/pLJzTz2T2b0Oi1jeo42VBZ/x2Bx3MC1opI5zS+RvmYhtg56pKHhlaab2G5GwCU6oGgkG/LHiJ2j
KHjKW7gsQteq0nnWaM2PvG51nq8LRJHIIeaJB1fpux2x5cPfQM9P7Hg3B6VsQkxlzhCiLAP9AgTW
2UcFjUuuPpYLBdKgV7OUjTWdwciFAk5HGdHD0lPgzMiRAaytE/vZTcxz76zqui6o2DuvckHF4Ijw
w6P9LdMp5AD2YQhmvBq2NcpGum1iyUpNrjvFNKEHb5rI5L7pnPTuGudmudHm0vHE5rGaVXOY6Y+1
XkUNZEU+VyLCJj4OyicnC4D766LKDPGic+l3WB4jd1IoPfv+sPq2R0/074xupFmJfWNr05OHlofK
qmCYNB2uI6J8z9gLuCZrNHI5U7rqCG2zl2I9WFP4YS6Nu+ct/ooGiSxsrWNYJhpB+MNzyzp6tP51
+wAK7tpicHwh8ZujXMIUMiVkCGqTGYK//64tASva8YJGyyk8J5JhzEEJw+jGEWWIM4KnMwoWabfd
Om0qdCVv+fIEY+En79exJisEKmYWQ0xCGx9JzotjzDxlsMqCzF/+Q9QMaRTGIBKoq2B0ssy1qrsf
ev4NR6VbShLc0m0YI2OKyciM6uS3jskGnw9mgM+Tm18h4QdwLUM924jlacmDkSelMjOcOXbIpZO3
ONb5o3lxCQuQfjd4EvNp0UmlmEa0pfKYELyqeZ9SjP3f26Xc97ktv5+pn6nfM0Tttm1GZcw/zcNn
0F+vKwvHNWTA2Bku9iwBISm7zxqUXHpf1nESpwmLxYO29lHgFpnkBaD6JtszKvi+MoOH/cRSmUFg
3aI/6EwEA4pU3jViWXdTvOlcZ+mJB4TXKh5FC15iN+KxpTmVgL/5njJH84gNL9zGgqJZR3D1yp5y
Oldvx3kFY1opbx8N6ItxPzJsjCDYK+4T3to7L9f2lorPZQ9ljNmrKvn8eFHo9FElHofI50jUDoF/
9UR4eO9pI6lhHmy03T4efoUchdFWZsu4hnb2JT57xyiUAtadd6r6KJpSqQV04XG/5EkxRBHmX9N1
t0+UmjG1EOGtHlqUkpP9Z1NrNoxPsJCxB2q1VfaoRYUhWIS6OGnICHqQZHeGCRim99xTelHO9oiL
R2y+EcsrMOYPD5RooyoE6w9jed/9oVIOXXi4dvP4j4iMQtavDJevulC4AMBGKef8qNSk5EOewa8Q
Xl9R4gK52SOvSdZ9FXRS7ZX7YDCCpcUdrBW7T2DvnivGCmvSLgJ0kdUT2/3OU8SUcbnc7IM0wvcj
eCumxkuXI27PjMwVQr0mZOwf+tarAM6yAFvN2yRVjcFTKIhnLvVFTJFk7yPV2KBVJlv1Ly5CajFB
/liSREWkmjTyuRqMJ7d5dp4iqGNB2klHa73MgoHftw4Oo/pHEbcX4u0a6DOECiTTkvqhcEoR0O6S
AOxwWwEtGFBIL+lJQ12RYY0EKqMC3XB15NB5WtO9pj5ttjQHevL+Kx/DwNCU6g+CYN0DrhAphJEi
5bFoOQVp8FM2KSRcdjYArmr3xICnnGjs2RylRNzyHKHG+TcQhgzWg0xVeXN42uc6P2VJGM+OrQhs
7DTSwL8gAgPWlGxFD+FQ3rJeTqFQ8bQ3yxNB0fcFJcbRdlKlFu7TLEbygli/4faZC5jRQ10RG9Uf
H328dikgbxEiL3tDOaYsdHxmRzdvp/fL24h47klcsIhDJs7GPtluXQ9d74LrDBVOzK4n7rZu6uV8
5ICCWKH4/GUT+PsvaTkWchR/0PideqjHq2Z6KfQte44HghHTevKjo7G4fvZjZxMZpRl7t92pXSmC
k6qiYluor7qjWPqdvoKCuCdcGxMsh6oX7W8HW+hVeE1F4PM4EEl9OPuTtJOI9VfRqhvQBTrIhqPQ
eOTTiuU1Rjg6BXK/IPS7kMcQzB203yY273qqe1S3u2inJufMLRZw+9u7I2ejpCTf+XC6wJ/MPRDP
VgNqOwWxqv5FD9Dz2Awp8PNvYHWIDoih/AV/1vTlQ/Dna/elKQnmwTYw5SImgc5/Yifxmj0yASud
1OAh1r0vvwfys7IIHtt8cioVz+TL81WAjIFh3FMg7d2fUIhg60jVivaUaGz+/U78q6KCX1V4Gy7N
JlatKh76j0qQHFyE1dWYtCs4Aj5HqLBXvsBqziUeEs77eKUNMqwOy96G4fI0MuWLNNf32xPKS6Ty
ycW5SECIl4UqEcn16IMVop+cXQ3eTvxMDjzQw6U/nSIxRxpdNyMQBlmiw53khihwPvkbmXGIMJrL
3/l7vcAJ5M2vgUlf4H0IqxJAxN+MZRPs9tpOby9Os3Q0kNCjKWUDelaW2ZK24UIzDB18swjozGXM
cI3WsEHjf1MUSngBxi2n+8brE56s1QRjpRbUT1bcNO6J+KY9KZ/H0sJx0yTnomsIbuQNwaixmzh2
5sKAeDGoNymxAudXJCwAzIeONWWhyQ8P7OJcCB0GxRwqLJ9W+c0EIWODFmwZd9frB5tyE8ebcClc
xxT1UA1moTLVXKHblV8O1iiVBdimRtBq2M7RljJ0Q2y9LHcLK1X8KxvPoI+OK8NPg7eDaEuL0+4k
BzcC6SRnVcO6URGcctXEhku5sSqjZDNzfH4mtQxkInHFulZiq1xhvCbZd9MHCNko3xgF3JBAP7Xd
63FjZa80wIC5syUYhJ62pyNhlPUfWcRogixCopoikabv7qUe4lyRCUgE0ESi5OJozn4i1av9MP8u
y3hMtWv43dwZqmf8Pd0VhH2+3nepBrkFvym4/TEq3WtF6KIHKa7oMIz/nG0aToShGoHcFNVInemL
12bf/gH44qcQAlcKDeiZVgw+pIMya8iBr/WB4ZPy3Kq0L+7wL/xYBih7N+rubtWcdj8IZrFe7sBW
TPWEn3Veh6dxF7DbB2wGBKNbuzsSWhzai95/8riRbDveuAd8YcPrb8VpaIA65hSd6yOdUs9gT2LI
M3CyCZaytlHpkx3UmGoB4vuY+CEVwtk5oFQH4yNdbX42w7GqS6TW4URlLDIxR6na6M+3wrZ2/0qd
kZ/wuKzP774VIanfzHImrfH3dAsnPNrdK22BQsb9i/w4orPDo8TwodaU+6H/RhDmlXcgOFTsyAxY
9NIvCGuyzBymbju7nznduUhSkjC+kjOypnuqNm/NwpN0R2Ey1upKkKypyRCC+APedW/jHeDNI/Ug
mIKUEupaSxkyV1WYkM4XBJnZ4LVwF/ARlUEn5bbNXQyJ3IVEzzyMwgmtBYPM9X7mpIy0AxsFhLup
eVezbF5YOFx4fk2qPtZOA/UE/cJT+6Kayg9Rgp/2JNRqUe3Vz7eQ/VAd+t2Yzz1Oigb/LpexvU/s
/cf7guyiZe9TVT3kP1ar6dhiYEF9EfbJFlhoATWafmu0XpsBMPVfF4SJMcX4VjNbgG1RTZvvVmb5
jaYff2T+2lZzOXvKA66R3twLnUAyNO5vVtLC2xPkKX8dF4FLiHkWvsyL6f9TBgXqt7MyHCrM41GA
pTDCbYFTNYa7x4ad4KtjUjFVhyx6uskBzfvXQPiLGOu8Zv8/EelG1b6YlmDTR/4ohbaRTmgBMLsa
kW3KACJzkcv9kh5QqzDIC9hDFlGR8Maf7mcwFzjbY7FRm0PFYXPXMzaKnQCNRrTKqZPPLfPa3n19
1QA2e36KstPkE3Vqi0o045MihYi7kWkw08er4UyFhMoOQe3NXRHGDW2XfAFRjMo4VIU4TMNVUIry
RKqRY97Yk0zvDrfGlazvuSK/yYVw8EbnyZGkZFMwz4dk+U2oLO7StN6IjUPjickP8/DX8qRxQl0g
zCpCrrlFjb+20aa+jXnLO+EFN7t1HvV7vYKjL6r9nBoHL0P86oyGQIK0V7N8pkkZaOFoSSHuyrOi
O1QtRnmPDPc/3WKx3dfFh2R1jr2XZMEXr1SwVEo9u7DHa4oRvrEiCUcFH3FOthUfeBEPTD+4gAWo
/b5onoBJujU8msug2Ntln942ZC2gbleHzQU3RhQpElp01rBozkLYLBlt9ClP3g73blTaLsijAjNc
8gEe/CEgGFE+wPEGf3ctTaZC6KzR3KQGQO0g9SM9ffzgfgCe+alFJaKeDQoVwm1NC8uLMtzgoxNa
5uWq4owUY2KkDNtTZFewF3dJCr4rV6ZSC2nsZQhUJ2NoGaJdoGsTyDimyipmwk6j9EgKZ8/iXqt5
xI8hRuvZQFx6WeG997shAe/a4CT7EWiKl6Fes1vLtsU4cocFsVacxr9nL5zaAvm7x74/WzzzJfty
KcIaXFHxNLjfJ/vx8joUpSQBc3uqqzDCdgrvJiRg5mYdo8nji1nWclsGJTXnDHkw/u++tjoUXDFK
Xjey2ipkdcxGspIFhbTf21/P32d6WQySDWk1hh3BBhiLD3gcEYKGV6Rf803g3FSm05TXjmKdDfYh
umsPgSuRkDPv7MAunxcIqihhFzb6hnrldaIlkYH7btxlthR/WQBC97WAWWJLQi9SwQhC71xVYCZ1
sUeenm9VhVmw8i0uOE3CR3ON5lvdrT1mBSEUI6LN44Noe26xOYOFmOcaOnATXnBeSxMqpNzx1j8y
JS7gpslkHnGna2KSTDE/zqXAq+hgmVwWTqp25SOiX1iyyM4JvZZ0VQ65sOyH8oypiZBlkZtc7csm
AlxYs17B0dXSM3FO3PhNY4Tdt4CEEqcu174EVWlS+rS9WVHXpJi8OkaaTwZZSB+appX50fX9617w
Qf/QrGhO8xoWeTljQkQroqMWqVbBLx0M3Dn9OWc/UXHXHYOhm2BoWgAr7OlpqUJDf6+mSt+cy3cA
vieTP1SfjzsTuOgvQkBz80PdvlEU+t3JjzG6ERRyazvitxgAy48ucONg9BrhS5YW2QOjzEXmMfV6
hcrPHsD0ZIZLoPZpwA8AyPgP4E+3w/4H52Oif61jQlTZfQnen85zMj5YQHTvZxq9IaJZ2+M3HJzO
vmVa11o74MK5mxpz3aStlnWgAtxWIDwmdf+SNAKU+4/2VJtcVLm+hnR4lnz71YwjCnM7f94gfOBr
7NDAVpBaOFS+JqqspizYA00ralRio/Bfxx9plKW1EX8fFmBTT0XcMED5C2/jkUlE6A4LQN6UPbe6
NjJqJm5H0D9yP2rXP5RhLHUF97Cf/LHjjMDPScN2if6w6CnC1TXemvF68gBUxrT71NhhVlzwXf+Q
zSr/9GkBwnjyQk5mw42du35JvjBpk5Fc1Rv2VROkNylTF3XBjI7gT6xqrEUysuHbSfhPhpKkuBYC
Yejvjel5g2m/j4wwtS/u5yCW3kpUTTzIfK7tGWPRKUQ+gmr7Tk6dPkhL7xIYvTBR6BF6YZ3x07lF
Sh36NQia0K9ZcfJeSFh0B7R+qucvSvDCaENh2WKMqaVVE5CFsr87x/bEqznuiAOqx7gXmvmlHmYS
Q82rpPvqh7wPsXoHMOS78rllpsVPSE0G9o7/TPoblfqgkk4GMKBkToJy7/A1k+k3RJ/ujY2CSLm3
AcuFxpZ7SQOLXv52R0c00MwAyrDac1bAbIkRIqCd+GbjA6K435m8ho0F+PkkE5iLHRHhJnAmUrQi
KUvBesxWrvrPbFCD/vjp3j1Pe4WfLwun/6YrLmQHHMZMFJBvEEaFGmzgOJsThbGv/8sVi1Pc7L1L
gzW4b6CDvStSSRcLav/ZRvcnBj5A9Cfk/JRP8hxU1XfBiklC7qRRbedzYdagYPjdFy5zWHiDBUs0
0/fzdNnnbSoMD83y/TORIoJpy6G5o6n9AoystHtb7+BgVmYd20x82FDYII3qbr7X7iqJP3nVFkA2
X+i4Ivu97GeB+sF7tUEoUIZLrBO/Bm2rcudr+ExQd2hY9HQgIID3m1x5oKQSytE+y8o27DSZkvBn
EgGOkbWblWmeXZoBdf070cc1VsHNfCZ2B3S57Ro2NRkjG7/4sz9DbBxqF7GnYh3xQPfRdaZAt2R3
+Ty25AG42K2kvGngIrJU+NsX8qYbKSFX5ZBi98/KhHVSPthL70uv658n6dpe1xg0n+HVPcCydBNs
Pc32TZ836dfQ2bCWctUtxo6E5AXJH8keiflgiPjfqdp24gwH2w1S0G69QeX2uKiqvyAR3GgK1/et
Fqz41lh7O8DoBS5P6F9NME9nL9Xr0WVCJf4uv58JIAkBfeNihckOdr9/ih+5vZnZtN1NkM4Rw449
EKb6TKmEOyKVeIrF4Cv492QcXydePs2xt6p3lj6Ndi8kE8jWfZCQyRRmiqzgFLQig4OYZ44uOlRS
QT5X/KOYa2bTG4ghT4YNL8jT3QWPFIEYherAMdvtHTfLEhOwT+6pyqaknOadq7xvbBNebIkH3yEB
R7eKpGg9AfHhDJFEZIQGSdiHa61F44ftofLJL6q2rXyS6xRMlOvgq61Tildw+lC8EbBkLjppuslf
8wlHttrRte0D6ZveuneWQTc6+GDMTSXp+OHSFlW83bOs9XvLWCzIfk14hEDbgDaV2kAz6WGjmidX
RXoe6PwFukG2kuYr89JUbpNrlN9wsf2CLNm5CRGZKeAqbFO44MSydItY56jFIDbfq5haC7nkeEsN
MeJgQkWw6CDIaU3+qHkmRvBnTpoWhJJkRJVT6kdjLdij8Dzeqm9MSSbbA+8dWmSbWloQ8E658UzN
M+ct3rim2h/2GB/JAYmKm31kInOZES3rThxvUQZJ4m7/WkiCjIQxJCqv7msOe3HeDRV2+Qde5nZY
F3gvhbg8GiFmzppTkJX0Suy7tmgSEfgklCcqxtsR16K9vk7vzl/QA3K+v9ZJ1zez/rWcR+fwJnUH
hX8dsiwgQm6Ez2khjep0TJJdnwwkW0u19JMeuLALhjkF/cdjpeEwerpGyfYHENV6ZDKkC6tCnh2T
r1sPWr0G6PPWjcmXPwGsGzxk3zdfLt2UFmsKWRwv68e9B81FPu1DmKj6PbPH7zxQuwYYz0OaZnrI
89ZjX/f/2jqWHr/EIM17lVSGPytMsQwsmfM+bQ1ETxbdA9CgigypmnnYfRoBFZhJrT8UqnAsWbjZ
6nqKlP5zJnK69v41uuZS6VZBcg5iaC+YRobYrpehZ1ltsd+g0JSeUZoyDLX+Lhus2QKnMYCsBUBe
7v/XUysJQsDgSLG9JPV2UWd77wuxVxMxVXDizx5pQ40IPoDGtS/Dx0ZtCyIASwZ+G2KGwDkIkUpf
9Th5pXYLjq2swW6+zpwsA9W6uUiaJUZ8nJ7rI7VpFF+GI2kAn6cJQ8RQV70poMPdjiI5gFheIB10
unPeaTHwl4OMFOKBodgzKRuNRbAq+AuALEMnTZuurp3jtWTED9fpllA1sEVlI447Mi9MgaB/JoXK
GwZxpyrM2DgkU2wnJEWCjVlKncn1pMPDPpLke2elh0GJuyHZceL7l/9u/8d3tyR9UC8yR4Jy7p27
8IjCidvyDbu/XVVC1tjWbwOgbD0pz2CVznTDnpjbgH29RjAzXCj+7OZOdsoOX1Da88thEwmkp9ZB
fc+66ekYsaa8O8asX1RLIeufKNbC/YCPYQeyo0u35XqxYw2kNLZhfwNkO5EPU82/TJMqi4/hrBl8
6sAMrxFQhyr/SodirDSNQp6aLwv2bb5AmIuN7stSCjJSJtZwSoUyLXGzqPBnTpU/9Dv4fgy+KfZR
1Ymmqx0cf1WGuqtqX7c5ZU/oSJIVUBXybbF1UMwht12DiKv6TuMas50Dhtg5mOzWxOWrSMolcLO1
NH6e/wPV2Dz1mBTQLUrzE/4AeBJnA0lRUmIlaJGfsKnSGWkdDagUsAIdeMDzSgK7UjVoqvIiGGYR
KGq1OR0w+eRQJAyAVpj4m9yR7f8av/4vEDTeZTv1bridNb9UXDhBZOSvS3bdwwapgkiHPIpMmryF
efiwIwIyNUTsWFMAACfeWbFjavnUHOAhnO1jOKFP4vC/l30c9Uj4kBBhY1I5YiAZPSdJ/U9g4FiB
H03bVYzx4yYUtrkAIrPT9QkRQ1Ba4tBQiJCgB/uCLfUJ+bYHfWnVpvp+NSlH4+Nw+wI2fAx9LIwf
5RPyY6nuxTqlSq/XqaCjAVgB68k7wz3LmvLxVq/qhLNrK8XsWpWLxGulKNN3DOqWLjwJAx3h0qOI
/Glhj11mXZ6DviJbIWURvNqHG5RPpLUVNrPGoidLJEGdWPJZQ5OYUauiTTWi7pqiAVFd9PJEs4FM
VrHxbif1MybQcpx9ql8RENh16xoMU222eL1Az5rbcWbf9CHRCjhLMe8i8aYsLjetHe4UtEFL64l1
00+inHyj7NcEFnZZuhPm6O/7emZJLUCatCdcfk7DcQU2CUatUh1xzmcqiPfULK6JyIQqJoqoxQQb
lbTyVdXVxOC7c+XZQjRZ2dpIaNOIQwY3brjWxuAzkJDxKjEx4R4TEy4dHTtOfQd413IRXMCKEI5f
C4i4fJ2dbahIPCcORNY4Fix7mfu3IXDXVfVRm52k2ZbEStPpGTmincrWl6p0droRmTPbkM6voMke
jygyLxg7PwLj2hNE4nvSGVwZ1iJbLDhxkZ47PMySFEbyj7KBaKMnDvnSiIcLo06dmdOJpmo3SI40
RW046Du2+sIbvk3fQ5UAJieG+YnZXQ6T47nH5qJga8C5UkduitHW31xf21/yV5O0dwL3PNw7vYY2
NXeK1vTGhPOKouQsf6lNJS92XiwZcKoX8EoQ45EqSmQF9uuc8mw68GnlaCNVXi3C/BEdP1I6yQXQ
x3QnXik13BKS+lJEgkwLv+ji6x2G3tWYPTCbPNu4qtigzFmubuBl8XQqGPNi94yIGotwPlD1Z//R
pLdmGt3cFa9ftxm/UHlHcnW/dwHp7gtJkolZ6D0MtesDqka74J7PeGXMaeDNFAyutjwykVV6Osx1
uuQQDM9TNaQt7aO4IINkkEAej7hK9zoqvxdXUQ4Qc9wzj296BBwor3fb51wjNgLPIG3YrUSd9MSx
FOZCu0QVgAPVlyXZjk53hD0U2B9wJxHJqKDlv5fveHdCSXLgP3zAPohOeB5NBNyQjwVp1xAKvKD9
zEoZIyLi6eO5aE/4tJU/BGQr0mQ+Q8OvfOYxdASVaqGM4hRS8VUhFSBfgUDLrVFiN0f4ww5JuIgc
oLX3KbpAtyqnjIp0mnkDqMRpsshTRrJcZYwjac/x5m7DO6Ng7hDGiXhOTmhweUOyQab5AusJa0R4
YwXOsEmIgrHXxzrGksK9IRVYYnBQ725T56ynj4li0W7QdN7mAVgPFlYZZOLjOxwuEoAcjH1m+x4X
mF7OcWNd2VJMbKqofgIgzPZmmvm/HPfJOFb73LOJoeCri+GvoMg8DbRaBVarC/0n0M0uXdKWcKhL
WSiAlSBhSkk+O6/PsKDiLUPgEz+EL9sh9wsUVT8EQAdjM52z6mDIF8NCe1fLjP9JPtG7js94s1Sf
3wzYg4V0dteiixvsqj1giK/qQqH6fGx7pTX6BGK13BLq5FPjCTkJcYPf9aMlzVx3SKhPegvrj9IQ
YXNbaUtUs6IbC8BEW04xrdAvtrpsGYlZoaTmbezqlQqBQM027NWq+3SWbXIcQFWAt1Ud+k1hf+md
gqnt10F5s7fvm5C6DkpU1BLBy6Va7zvPxosez1bq+q4OIphHWS9uOWdev5Lx9sEM/KfVMUo8S5EM
GjmOtApnAMG/bfTDCyB5qXdaum+l7P05ojlPNWwb/SD8C4nOJnfYT0adMxcSkthNQxdwYhSBvxB1
SAz0WvmKAkHz0o2Su4jPMhWGDlsTp0VbjCfsC3MnaJ+OyKwsK5wHeoNSSSEleNJWdALtmSvF5iHb
uaZzv0qMuEULiMFr4oRR6NWDG/d4mpf2gzv3ayaSRnUpAuw6mRc/0fqpPmeJcuBS9a8sVOpXJ8uN
ECEmvMP+8eSXYCpFWswqqxHj8WAs2lsfASXJpSqpHZNGbSnHqICHC0ogfj/7CI+Db4uUdeBuuMUK
VvzrqE5h2pH/vF22ulJZomBLX1PyZTr19aAN48cG3CK9Rdauoz8u4Z8hFOOSVm5NhX2FrV2D5mkO
Ejw/iVfjYofMBUt5SzTSYvFygF6m8XF3E5LM5sPupBhnx0evkj70dSzVpi8nfRlHzSw0102jpGIr
dF4CKIAuvP2Fh4ekudV/C56keVU3LUmjU7GACZ0YiXBbiIhLqpfXI+bMI8w1r5ALZQ+er0CEgRsU
z3sXOXGyOVRJ8AKDCzXtmE/Jq0IMdBFlcZbZwI58ZjxStni21fM5Q5d4rCID/h6derlkuJkYe/pI
+B85svrUPyPLYLa9w9JBM1Doc34kUnNf9by0DYjIVTj9boLXWeSvhwTMW389ghOcAdmLaZnsuoC7
laJp+hFGO5MpSuzhaFj6+zTUtStLhZFsxvocgRo0wiaIeGG1sM9Oi2mn/gI5dO2r7zcV2QVBvOV4
BkeUBI8X4mrxwqE5vXxqD4zekhMI5/c37gZHM/DEwK3XovsiOzU3rIQCUyVIp5GOxS4sSLoRdw2F
WyN/SxNy0hiv6GPUurDjZ7oWHv6K/r0cwEc8Fs45EKkLcKMj/10l4SXTrLRg2dQamP09kJRY3dJ1
d1WY423fLdtfQDMK2qbRyforhNCr9UqUcfZq46pLRDO2DyWUoE2bLzSTHpWMjglNFFdfkCwIY52H
qNCQMmRxIoxHnDD+jzZpO0szqVIVWRlgoqbGQcA8UDw7IzvGF415QxcNVa9a/HUBhIS9vtDaSMWH
eKe9Nql1OBuCLqdaNbeD/+L+PAy3RxeIh53PFHJSAA8Qg0jNTmNsDr3tj+uJYX0ZuwXWITHa0P6G
XDCE+HUvUaKs6iNpuOqbmFX89WCtjo8dsYXH+SW0uLVxZokyIq8Tdqv4anhCeH49y6bNB6rhx8ku
11mFfYn2Wrqws6gOUbbEcQ/UIbFHwchr9AbJHTaXxPK/z7cRSWjss4QYNHK03MnuYhgh0pk/fokZ
8HPIngpl3+EJiRh8LgmXBsV7lor/KBi0uNhNqfnRW9a4XGFs5SS+KN7fUbmNp+Rz5F2wEzX62vNt
AqAoPBHP34msEAurvsUYVLMycYMBqlQHal6zFWp2DlC2ZKylQVZlKfPTiovNeiHpDhvsgipizkP2
Jd/fxJTJf8YKfjRYZA2syDJeC916lvJwVu09q6qYRFWnBN5Qp/539kGrPYAPd9mrUsLoYirPenrz
L1RGgl42OmUBTaVR+Iu+KaTilSZ9IfPnnLs24kZ6xc9XgmNsu4tV15hQcT/2auooDaPMrum5R2nz
5216R+/WC3JyR4xlGWTf+lgTPbRpR+UqX+cl7GjzMHHXs7dEpiEF5XbPDC83+3zldKHdFkd5ClQp
PLCGQdjejj5E3DFMGFTp+m/rh3PZMOOK0G2Z814Cx6zdTCO3YGTCGZ6CemlOc+E78ZAsxW0p2n2h
NNcDVgp0tul59N1scxpgwiCLQVQCOgATOGdMdBGNjDe5T7e3hv5fzu4vUoDYY8rOxICMbqxmC0OC
J3Jyq6JZc8nc8Wmh6V8e/yu7Hs6qa7IAk7WavFq/dePfazHMHIXk4BgiLffCb3zQy+DWjpylui59
zE8piIPcsXoPYWmbW65Ixi3YuiZmka81mCbzOHftmHXIjJvBDorK0rkW/PeotOoAH3RuWRlzDW5n
TceObJdjvdlgfutuaUxL9lx13/0vmnnWko9zy6ySRuCTvyuZHOjBddt0kRot1+qTAeaM6VaAQUYB
l7/A4twoqvfPmHwB9u3QLFrYJ4br48M3VS4jXHK4ziIFcoP4AThcwozlXZv5klba74EQ2NGd1ZUL
qC+i1slv+5Q+UrIFNHj3TH6+z/6Xff3kWXC87g4vbif84gclsQ5q5MANN1yOpukzNLhhjwAHh76p
v8rtUUFRhLjbRa9eiTFNceoag8v0v3svp4LDVBwblSPVWQg4ADxkcEtZYb5aWPv/NyPpV9ICW50e
j/jen4TdR7B9kXFCw8IsPDHDMvB6vASxZ7F161a3kPmHhnXi4tHPMDHGOaR5uyE/BudgYw61MUJG
Wlerd1vclr722KVZ5zBmDBac/PBE2k13ZecyzAgox2y2dQt3KgZJ7CgafnE+G0Gyqpeaz3nJ7DAd
mo7NY5LlVcbhF4c9elOcKwCpF1qnVahI7thax+51r4YZWGas0oZjhjejd4xlDH4e6Z1B0OZ/gShj
pBA9XVZkczPTGIZsLo7gALHLtRp1nqFJw2y38YkS5OXdtc+IMcAxVGFvNHnf98q3viCUlQaawxYx
apmXzEr4L+2ezOgSr1WF0OP0WiGJDRvUib2OSxE68u3kvqmA2uO/Yrj8YsHr0fbkUWfpyXTlFcJv
YQnYBs6K/kb4iz6IiKOaXL0G1ktWpB9wW9m7fdRjpUHMc9KtfBbSHF/wYUDG9QlECZH4TVFqdTBm
oyJPF043GtdjQ3oTmo2fqvty6hKeY17TFbj9GN9J24o1e7Fq82zpxaDal6NKUjqu9F2ILW6blnHY
igi91hM9A0RAvc5lBR90SGnUsjad4wHLvkq6G/1G6CJVM89hyPJhP6Wu22WxACuCGgLip870iFIP
sFhPd2x1j/AVPtKjN/KnBmHRnVilC4t7zznEoRQ8587mAo//Vjfm01Ni1FrtaOhJkggC36C0ud+l
x0jebFQYxyksMBNkCamm2l6mVEUzxf/Xa69U1uBV+7oSV7PMBOgL51Ay4st+lUXbbenKDUmAacNM
q++FLFcqSwdHez99dAx9SI8gIkURKKpInH1ZrCB8E9PsnJkNZSGXXOpr64kDnZ+dMN5o+2exoB4M
04e95UpvNQmPctOwrOcTi8Wg3T40Wu7cqInrGI8b8UHhmgvUtxOuJh6VvV3yjWcqOhd/bPuaKseJ
IMXePGiJhg5iZbTix/CU6q0YSRXJqG4RwKhGonV34m1PWPjupxnEkBt2fG6WsHPQU/3sC+xP3YvR
9X1eoaCjQC7s6mrAeiRXjO9hXEf6hRT47v5BLD/yIG7x3Jx77KItgeFeIS65mLcJ7rNKEN1AhGno
hU2lex2h5mhqi8w0BSQakfuD8zW4qiYPO4c6FQj4PNPFRUtMxjhPRNEbOxJMVPFmn207cO8X8SHr
cqXanxqSrCo17YRV8hEC/FdtmXOzeXAQYV7S7JWu0UNaxep2RkZgA3p5N+QKV3w/JjRGfPr5yOJf
oJQWgGL1B16P529/+JO24erHwhuE2CE0OGAPwusyCfHxQZdkFsS90iXHF7jf8mueeWIESP5tAgtN
eIWx8KWFrXRIzmJhfyz9uVLHUgAGxv1XysI/SZ7h5Xnx766YmxUDIDH7DTbjEc6cmd09I28tJRtw
QiCgLUENeg/3rd+X2UqWxoD7dDQVR0UA+RDkpdnVbT8/vp49YHz8UXOOhLWFMH7FNjQDUhkPn5j0
FKSrugvFyzrJ+E5eW9UlDT88BZ8jHF+21eXTqhOBxjRSJvwwB1/i1WylYgkVN1JCMxZc3VO8/Tmc
NFs8RSO/p6SNU2Mgg/kqy4xgY2P9FZWM8jVzJMOgUFWSzP9CB4aUyHhRHCe2JrUziIA05T151uRB
MImgbyUBMM/cUn3z352mS63yFQYeqmz1fPpfTbZtDh50QdvO27yXerEr8GL8KuMv2fr/9MHbrxWM
j5sTnm2MYnVwyj8IOqltXWfaVpjOgNO+QtruZIHJ1wngPq6NnmJ2txU+lj5Gm0PVTwsQQ2mcBCV1
QHwEzVXsHSOCRII+41UX33aorYGcGaLCiMDXhxuAC18G3c4rYfwulHIHZ2YtstjtDWIN3a4A8EqW
Cn4hsWQENaQVOjxmCU5DRVY9438PBGONkglGrq8Fqu9f3oTAdok2fbgXBrOOED6mgDxX6zxuEzm7
dYyVF1jQjlbT31Hx7ISyWzPXUKlaNxCFhBgjxF0tqaCfH4oQuS9VZDHUGwqNALKZsKKrI6Zrisvf
vISbG224c5yYQgGHrrRCfH9OaOlyXLC90OrjVFNJXeZzF5RV+s3sWEtMBT5vhGmB3Ll9MNYQIL5m
mo1Aikq1fh6qnlF4A9zyU2Dz8UInrrDe+5CjNYAXRO8Zj73rai+EHvD85FZPb/IQ5p7yu1sFkn22
fux32fYfwtcy5wFVd9GlLzah/htq093jFYPG3dXNHYy834G0tt++dX6BHulh3kqiXfMZbWZfvYbW
kXtZm2063oTOatRNwk14w7kKLrj9eXCAyzxp2BkpcM8CK0r1EKv4+7FTqtusF0/1zoLsQ7qxn387
fRFGaQXpnRbVwRZRP+9I46M35jBXxSSnnlDX6Go+r2/6HKvIjo3TrkVcTvfYyPX33PANX1Fbwb4b
85NDRsvX5uwFdKTmJgJdl37D45BlRKtxK5OlQ8dHt9mnfrIaKgat7j1OVKe1moxT0o3CZyq6EVs9
MDu88ukfZZugYV1FKxCVzebLDSwzZofLVkFIqDwn0ycyVbSdkwmgtPZ9s5aXpiM8X5trX6FYYcn8
jaNDm5g3LXBegh3rNwdwhmijNqM6BvoQTpv6qwISAuObV6JoVVZl7+yC/t4eqRdGfKFKLBlpOxE/
5X/JnmwPcd5gjheP9HEDumKj18ZOAeamiFU+iaPiwoiI38geMVhR2dZT1pzJC5tjUkScc5lHgoHQ
H2K0YIEItbH7yc7Jc/b2FanBJpmFMXdT4VSdGnbDdr0GZHGhKfRuWmnM9dPGy9DuQiUomWFXHcve
9miBawPA4yI9o+mT4dSSLceAoESMQZyOUzT8UgCF3HgIQCQJX+lmkzJLIk8jPhymTd3lOgERrfYL
DndirYN6kgJjIy8T3d4wy35drZdXZRB3wsQETZTII9zz0pI+OL30cCDgycuzNpCHhfftg/WTgk2e
qdVM5W7fmNWxU/Q9GkZ55QAApkMY0ilJolfKGdQwPoTBA6TxkDkQjR4ieKhokCzsuxjvhOsEU1x5
1MkohhmQEYgvKh2pOjLiP3sw/FhBlIWRMD97Z6uKQt+yOWUAOTVSI9nibZ4VkL41k90Dj3i4lF7D
zyTcsAFdOkBZeM9CnQ7xljQmjNzGio39VsNFGYxVYo6DZlFHavwXfCrqnL2mJmmh02p7iIdpflwq
DWw7qyhlYaeqxKtg/XhPnppDhgNJNOCnHa+JtqknqNlf1wPj2Rocn43oX9qVGSLnrf341LJgLD92
RKVs3wy6mIXBgb9/1PVpiSrrWB8ZkZxjTtx3SA5NHA5SOZBcNBcs7dG+pGgIydVrl6DfijGz48FD
7+ZTgBpQ3BrMLJxisIZ0ZI2FQT3dRjsVLBEEoYVMHUZ85eAYnxXFVQcYZdOrMITDlLFPKCf0TzHB
3gKCXkqawvaJD1Ep0Eq7Dqwjwf4eLLCX1T0T0lOtkuWHMSKfVpfTGPAnVyPudFEGFQuXgLqjVAw8
BZeW8JI7Ob7/RR5iwozbLSfQTvPvYTxKE9YgefVo5j1GEV7fIqaA24KVpWZzyHue16kDs80jXjeQ
dg6j8YX+OEd44n0NZby63GqJDssE0g6iqt1h3ygObRJkr7LVldHtwaIhwUOGq0IRCqI1xUNHyzV1
r+3tKXUpvpsc4ZXJtD3ldNufDomojGGW5OrYpgnkH/EV/Xl0hiD/1kCmMBGQ2sSYQ4uQPDabrOC9
h5G3+qXO5dvfNacaA7fGTyE4Yex7wYRXhNHEVQBTklEUIHIOM5Trv5FMNI0nP06ddU7n6JjoENtA
0qCRxZtrxNF9k6m7Dahp5w4gj3/NYT2s62GxxdClFyW87DWVItuPQSMlienJLZWI8gliDYkZcNUB
zd6F2gSGx7OMwwTYs0AYBIfopphwf8MDTEQAxYjlMfNfUsqnQKHspeOECEwmtSSf5gVK6+33+8zS
/WkELgeQzACYMxIGOfyCY+YzV8XRO4eMVOaZxQcnC9Y5wvjyZPMntkcU2XCY+5l22ow/DgCqzQSb
JgNf5Hi33GoU86lyqqXsjiycCMqyQobMCwrKjb7b1yvb4kJmxuSnrdBNfeJ6tE471OHiyqArzntF
ANBscsNPuq1WXbbcZTzFb3R2qethSeJPpQ29MVYY2BG1FipiBqL0/b9CYcYs3WBFic+IH8+mp60K
zY7K4AdG7LaajxWO71VnpHnbRPevh0s7YdprANcSl5OmBbatSlASMXZFmXwlkzo1yZcMQGL5sTso
tdrXdspfDFwVAxfzIw/hQUGzWpQiIyHDmS6BQWdRAy9YMve0gWHncPYGs5kOirpBa4FvooucRNYy
mPe3+UlpEptkXpV3JFTbIjq5Mt26FrzUSYSEcHn/228fe+4gBBsOuQb6g0YCDmWVBgwX9VPNvUlK
Cx/1gzKvW+Tq4pPPFQNHtAIdHNNCoUNM/C091RLWIA0hX7FRURYj3ZIffUNBMEXidp7/kh4ZFNRO
CEQBKlM86ehdlh78w8E3dte/N3Uf+c1XDlPXaUkdjUgtXJ0/JS9gqv0CSg07OTlvl7nDP39GF1gF
433thIbDFcrO42ISf1+uj9iGIFaKBJKf40tFSB7E7AuPCscw5s1iK3dS1S/CuAwYWhxhXkOVOm7e
Tzre99yMceFfasIOhXzS66/TTtcrrUCXJyhcaEh0+aeQ10rmJ9w9bHoS0YPlQpnRkbivkVvxYNA1
4CedZdqehh0JPa7ScBBKFtd8tg4bO1T1oC7mn1m/1JK9ndgprnMmOCFD7w2LYD/HwZUcGJM3r3W3
qE+k36vNlfLLEOoqyfMhhsgINPUhA73XJvpaYgWGju9o1teA/FzSSL9J3doArJ8XX6PsGn1/AHwL
3Y+YnFuP9kkglPt7loC+2XrTzKI8nnay1ltrnJcUIFB3e7Qf71w9IQ0Co7EeEeqa0gQpT0YjGKgp
zgiwC55b4Yrmw5dmgidhX1ILTDhf2gja5H722M0B58qOfP04FX09p9htXqlCYHDnbXBCMGeahtEC
6i+U9Oq0fCIz1ykVUvd6GhO86nUbQYwGvrV6RTW7RcTSbyg/mtIwDs+dwaOG4jBtDrMi/fDdY/mL
Nuz6smIWKCHvo+EUo508pAF59NeRnUrC3BturbwwmmRHhIFUFtAqnkqkAPjUJR4sh7rG5ktsePSc
0a11MpTf7a8CB+8OMe6m6ko5RMJ9Y80EhpkJ5ko1C2R4v4PTbYbnk62pN1NlIBXFdJP15IhxGJvA
KT9YjYxDx83CJeVmWA/doySZ6G21WFM5AVsx6479zKPK+cR8tTAKZPQAKKY7kwFXQt8zbyj3u8X3
k/cvbNHOSO383XvJEduDDSIzG2GPCxbLk6dKE82CRfFzrHcYxR/ekd6kUqXmldwcJoFCzw4RyPvn
C2n/f784yn4vc0P2V7lZuLxSuY0gqi6tj1M7Ja7ZaiZjjhXoWtXopvhgUfvgLA4t38jCi9nyKzrE
HXJwr+q3sQOHY8s37JZb/luxifzzk9GVtDX2kbcHFw2QGOWX1tNLe8cA5Ge182XRGVDipJb96/Jj
omko6iFV0zW6zaQQ38CJQfzSeloIEEvnJXVPsXHge5A3hvGIywGJ/g/buyfYw0MV7t9fCx8mztq4
McSCoV7bPUfL3+TWzBQL/rwzbfYL1w8HAWnRbEhTFHSMTsAvgmxpKqg2ENlq3kOb4LqEpgGmbZSF
kSx7zzvtkvkFDLKMQQ/VDUJmaQR33okna2azmSZq0FfbwN1Oa2lJzwJJoL79RMndHDZx08d2Fdye
hf8Xl1F2gK5fUjL+mxkhultIqjX6VXOs/qMwvQXBuADNhFDzR1E6PBLX+jgo+kNeAIdnCb4LbvSM
Hjc5RwO+R2dF5u2YGXRa9bG5TN/jKVStYqdtaFrV8Qit/zhND8Pc0OD8IPaabdR8vLx82CGpayki
kIpf5Cg4ZYjO2JRAghItGFC/qeIEq3H4Z7v3T0yHm26RrxbZlpqWbOFEqBPxTI5zIK/9QpOzjnMM
yLvWhc6/GLgsvKVQp8x1ZkupK8ZKnu6APaMlCZACiVH84S6LrhtDrPVtIOkQFlRQG7vzw+87MS/d
WZhee8fSrf8LMmpUdyBowA9aH2cSD8HmW1Tk52iJBxFY9mH7rO4Tb19+pzEyFE82P+qIVOVXlcIS
zt4oH7Y/O1WZu7JhbBs4SZf0K+gKXfTsLUVM+3jArhsu5fN7qpPXyXcD3PxkMbHnhxU0PN4wu+Pm
FrE4c1KtZzivjIOrzURF9lTDPl/Hby6sJ/ng14W0E2/b5kv3H4osv4Y4d9a6fZo1EeFvAXaI5JuW
bS0HHWABkHda7RuJsnGUk0Xnw6dqmo8SBNIF6UNf5gFtraxn1oJqYImW8b2JaSVL8B/lTm8rfLtS
LIjE0csjMh4Pfg7ntVGCsPvR/CNyxLqCoYF5dWJfUF2t2fu1hDjgOxUEKzKr6ZFhpyesSIgivOEZ
jK8EuE7vZwvQ1MQSI4spB+FDmv5ojbpE/Vtzia9hnu8/x3+4xhGp47U733gvO2c4wFyDYD0sojBN
u4hpTMUbthI8ooK3YbGM1KptQf22uMCw9+NOsybJjCvP5OY4xJRt3kBk7uHVSJSWQsXZm1EoKus0
wfH10+XAlzCgaXm1kJ3Ztjj5Xdv15DHmYPDt3qCtongnX6Sc+GwP+3WpwpEUvZH0ceS/3/+4pIQZ
rbUe9wzK2quP+C/IW91UkY40OZKVo8hwjCosHSi5wA2UMFfz2hrjgNF/K712jMszWGBw+S15khRF
tBBHJ2Al3mBJ9QTmwzqaKh0JjTUCV9SqziRzFpJDcHHlyNH+Vu12xr0V9QIlDYVqEbOTGYhPJAN3
ZY94rO43bATYjIuDyw1mXTy2cxso7QhhG4En4btxSp3PeQMTB+3EfbJsCFfigFomWX7UPLG1M6FO
ky6cg/VG3WYAGbn+vUJDIEmwkvAMePnejFmRFkJhyhkiYTHJ3R52zP1KZhWZBhqECpx5cEnnZIME
lgPI9z0MoSRTBAmlJouAYU+ccOsF1LMtxBvx/ySHwrP4kPp8Tcj/4q3agPQvvl+S8+CtpMfeRktm
HuOU+lUIucwbCqdRDdOwTXUvL39eb4sHwX00LGcIPBY+Zqz4JlrP5Im3ElxcIt0xgCnlqxeow6K4
POl/413o4iKm+24O4Y5BaRNpucOG5fs8ZMG6RYV0A6hcBQ3KS8meq/Hara5BIGo6mz14YIWu7xpM
6XVK2hV59JTNOyLzsjfWDnFghZrMK+86QlktNAgfuV6ADvmMy6Et8Su2QAbhVYfklMLBCnhykc3G
v0mJUZrOOrNVOKIZJbh+xRHH7H7xwvlhN748kVMNsWeRGTSAMgtkkkh1jOpp3iIn8Uqw6j4wwzcj
fxnmv+QbDTXwd0PLaQJ247z0OIWGR9MtIZc7KzHfIy9vSrbXJHp+rpwjVGYW+ePjd2jdFmMqIOZo
jmBMjtT9ugwy2gDPxT6EOaOtTpZeUBXWX0xxhGGNoqylXA+7i5Hxce/fRuVmBJBYQi0q4QM4YFXw
lVrf2iI/OD2700rOH0uiN1pUMsSX8tHL7PnfIbmq/4JZ9XAEEQbGSveYz4xhpPNnlRutwuV34Ilh
9v8YDVzi1Txs+PzJ3KuPiZAAJAG0raaQSniQGrXlhUIgY7GhSAGWKEpiHxw3FcF96i4I61K/9gbP
6a9XYUrINFwg6MGb7orDwm0X2RGZJkOyXzyqfIN59fCijRHuf/YpBMUI6COLZiPjvVt90lntehK4
fq0+Hzbnx0VDo6rKoSWKgl7OQnnNQ+6yCW0V3CUoC1WhH6AgBvi1gc/xE0z++6kwxVZKXdbv0dY8
tf4D5G9YTxvyG7W9V5LPYpoJTuB1CYigyPlYsJqFlPK8Y6id2g4Il9E5dKmEBvKBM0mrBbb5aL+V
UwgseRnHb/gWZv23C4W/VxvH0xPVdPSvwMgddaPpTkHns/RtLUf31iG6LbK8uYVPDoQI3vplexsQ
ME4UK5SmOjvrc5jy8+oDpcvT4Vrwh5vcFr0JuZFf5x0MJIXslxGLh4TeJmA6p4nf5TMRwyhWOMqD
uJEKjjo+uB6zhRlQIf+8DT5rCN1puGyRaWlJz7thtk87lirkZV317LHZahoq6YqUvVh46PoQSUKJ
3TN0wmDC/ABR98zASVHnuBeYq55/1j4rK7UiqWs5i5sClp1VoyOXWNe08kxGq/fUs5vAkvV5OBST
iChvHJNy4VGBU4Z90RyotmXNHG7OFyautbnJAoraKxg39P+shHf9BJ2RjOjm22HPnvYOzrix8xMd
r0kwTgnWo0gkZxgSfoHyBx5EHx4rVao/YsBqziLOVNy7+ZXzRjGw6I6++SK7+6hkIea4+0o0LfBM
Uw6SdQNYUCU2i/iI+gy071JO/ipojB0wSiDswuFphQYP8F6JBP4MZ7oAO0YtjrXD715XsZ/ZHQ87
ZIOC+oygDCzKselQdv+kKEU5zenKv4+/6PoGa4ct4QWgCg1IjQF/lcbxNYuGB1k+BVrIxNeITYt1
Mf/rwFmCMFXs8QDAZYvZclG4i6SdHpAJkHKB03Z680YhTtk8/4PahdbDtG3BJIWsImTJ1N6iKKa3
ekTTEG3nJNEbhYn8w3DJ9jUkFBnFcO66z3cpo/DC1IXscczH7ILnVopg9TtV7jtfhTlZkcrzW3Uc
5tbA/phX4Y6wNBvdhBKDANabMc0uUjsIexwfy+pXc0qBHVJOk2lf7gFiXETZ/m9v+N7okBdvTu7m
ofxmAKATtoBACcMnNo2UJrfz2GBSxpjVqvxRZthe6en6pKWjvQxT0P81/u06BMzf6UNQuYaEwgt6
27pB7hDT0vt6S7DoU4vI8YtQfAkJddmMgad13AW6YjfOLbQL6AmK4cPRPelT1UVQ+ajjafwLCBnR
tvmJl0Jl8B3Z6NJ8VMI1Sobie2whPMYvYemen/nDsNVzUZ35/BzTKIpjOHPRLyrOHT9agTdhO7mF
LkGYjHlw7395+6hQUlqcnGmdeVASRsmOCoVL3OUAr4cT7COcncC4tfFddc+V9bGpSgZ2qQ98T5FK
yFBMEYWPqy4A6OEdQSKoe3NWaq/rQukhVh7EMXxg6V+hYbMA/t+f5roQcNiTw4zoClRPQW8d9xI2
D7+sxelL0ZSQZMiraNYRsA2oJOBKeiwEDiJeVUc+xCZJWTblS8b0qZWkD4sk+iVPaUkLvI8mlQzk
QgsaTeeH6MMuW0WI920kz6mKXK/3vEZ917c7Fr+akpxFpcpfZDGoftQtA8bUiSuldtS9biExn61A
7aVqjrMF1vp8G6oHRKfB257HWsLKrjIoXk6viNVgc7GyTrbJuvw3coQXdcUyUWosBKXcZiooiSFO
XcUorjzVnsAM3MYXISFeip/1oCg2nJNnyZTMNMEvrbS5x0IAWYQDtVJtT7cyPpjzw7miUBEIbP7b
tH9cHmS7IabUtBuA4fskfmtvU5LUzjzylP3Xel5xm7JWb2Kk0rfoYIUzpb/RGX3hLyUxnjRz8QTB
12Dn9kJ5mlXox6RPi0za88WGDYlnllnoWGKWTElLlAijYxG8MxwfvrTqQvfQFPcn/BmlDlmKWD6j
W71wtMxKZZzDJXj8JFfxzTQgHTNAt1dyNKJspfApahg71ZZlshTEm0DCI93t7X3hqQXpxciv1B7Z
BBiZsLl4ilykx1uwRDc4SGkZTaa2GMOK7pyoFiHd0jGL35zDNF9ayOmduzDKC2VGh2A+hw/difNr
UGm9J1Cy8hfRT3eTN1iWbKrr3XDcsNnb2nKunqPXgO9O95D5A9bcLyGPk8Pe9Q2hIaC+/mNyUSVC
qGJ7pnnYkAaZYfrCXstO40xHGej5xZckBu3bGHYUMWXuyP+ARH6CojcW4UUJmQuo1NUqTz7e8E4n
HK/fz1Es8AILj9+Bm8q1ZlIAy2XJ+1Wv5uD5bQxGjzKekgunaxhMpIzd00xVtUYYnsR4TLxaR+2M
m4W0pDtT/++yTPCpDLmiD9jK3tjjy0PaO2KCbsiGkMT2oaOHGOImUodmzI+U6K6hmZpO86AQmmSK
F6q1csfCNZ0iLFvIQaSalEVyEilOSAfV6e+c12KyE6jbYDILI785Gfne89WzK9Hun01sK0CZsrOM
8t02/VYol33sUHehtM9s57tuI9mBOy1650i2CsyEnn9CgyZnpGC9RTbznB/+dFzJs9sb6VINwSk8
44tDwb9vB4lPoV6TJ5dkaFNg03nQRrXzh3zNyBZvsOagH+Cd6i+XcJMegDNjGKLg6rYCJoiB7D9W
AECCiPd6PAOLlgKr7n9Xz/4dYmcHBUHo5NKl1nRpZtwtnaBoL8Gsnbv68zpIa41X1QXTbSJZpeZs
yZJB5zxaKK6WoBYQynpLFrnWxgYW/oTTQyGlBhuerRo9pGIHxZTdKQE1MvR7g0v7KcHQyd2VW/y6
pqlq8YU1gdhgUvJqwaeFT1AUV2BSs7EQvlixswmp00hFf4LK7b1/FrU4JAc26v05G132lZA2PfXD
bmzt16jakq2ppBoyFTcB9LKLASipWebLxysTPoF95QtamtCLH8W5vRo/zDAz6XcMhrMx9FhjS2DG
hgi6RvMxsZbtSOXGJRgOHC/TRUx6GF10lUmoxUYAsYCkHM2lqWwUz7AAbaML/kKLM1PGov6LuDy+
ZxKw90i9Ws/gjSlZDHnOEt2S6Le7zj+exuA3VRj/2x0MTc5mlpfbttFp2Lv+5WQ9RI750/eLXjC/
HiHX72Y20UpZR7bDk4tgxj3Npnc3tKlAHmHm1qdFAyz4tTEXiqV6uwfX+KJQxiHLGxNIhg7104Pi
NEQVfd6wnmr8vGlRI8uaOCuvJphRWPTUaK7AcHfZ6faOK/lXVgyU613ecgIABaguivwzxRsr76gx
1kNzdUJz+5w8OmNpdqDxIS6m2zAlKY6VAu9c/jnous5RE6praoMoYyMXATzD/ifd+ZubDSHsTE0p
AKDCWoTQLAfh2ZQuRxByVzfkCwvH284+v+7k186KGwHd7Fsvy8C2d17rccU+4BpzenroftgDO6sl
UiAq60tk+rQ/yAVUsJ24U2J/JrVy4xqaDdqbT/KU4s5e5ebU/DPNeY26e0BVxr1vl/QitojD7J5J
tOne8PcecKJra8X/1c1/PCjZKvcW8cpVKg/X5d9aA6o8WzF90WjT06ewWVlwkwZymiQmEi8sXeBA
q3TJGMdS0w5ExZgjWOHGxEU2F21Gy5WrdXqjIwkCvaIr4xK+iXi9R2rDLyM6+iEArZGZMZnQzyKU
RPmQI0FlJuCjjQUdNv3OTTtrPnBltP3bKuuXeyMj4w8kOWZ3zlUatZ+wWTUYiex/FctoqpTv3xjM
zgJbIAK4C+bkt80/nf1scZicmatM34JoXhSyYo3cX9ag6zZqRMJ4Zw87jOUEb2ddwstETeHGfL5M
lPf6USvrSe51OxYsi2UdOKJqFkVegem8YT4OGDYEgt4RFq0c8amVD2zuotXf8K0jrjX0wOWSYwY+
VeWa000mmxRlUh1nhD2+HtQkz4w8nAGzhR6vURzGchc4ZFadyF3a2IMVWQWBmz7DwYxZOAHIKcGB
hGm/11GXJxdB5WmS5XdIlDFXIxcXwGCzYFQ3bHwy2Jsm4yttv7z/GHj+fXpBXYiIxiUMCdJcDeuk
EYHLm5fUz4uglp0LcRvo7hbesDZbwOW4YC6TUfaG++w1bcBeNajXFOYtR3bzCRV835SLsQxIuiHA
OjrUg+b6Vzs5oJoLnoRyGF862LrAES+v2ndi/eGfODtRk84q6PFiicrjtmJMW5ix7Pyf0eO2mgqk
kaYO12/JAUNKoT8mranBpc+jl6j/XS9bOoRudGe+1t1nYpGSh9VWhpMKMXH1cWoGVjhykcyC1tvY
WB0SBqh2uB+GtZacoo5vCYRe4/URLsrx8dq0ivj1G+zS8E4Vs78aPIBvjAaLjDkm5GeOzW14AFFq
IHX3Lf8gKi+3SqCQ9PAOazKSmF4IEbo6OqcBSX0162NQoT+iT5MwhIEw2M3M5NMV2ggEExvcx/5f
TRkYE8o=
`protect end_protected
